module BR(instruction, state, controlWord, nextState, K);
	input [31:0] instruction;
	input [1:0] state;
	
	output [28:0] controlWord;
	output [1:0] nextState;
	output [63:0] K;
	
	// SA = Rn, SB = Rm
	
	wire [1:0] Psel, Dsel;
	wire [4:0] DA, SA, SB, Fsel;
	wire regW, ramW, Bsel, PCsel, SL;
	
	assign Psel = 2'b11; //PC <- PC + in * 4
	assign DA = 5'b00000; //THIS IS A DON'T CARE
	assign SA = instruction[9:5];
	assign SB = 5'b00000; //THIS IS A DON'T CARE
	assign regW = 1'b0; //Do not write to register
	assign ramW = 1'b0; //Do not write to ram
	assign Bsel = 1'b0; //Pass B to ALU
	assign Fsel = 5'b00000; //THIS IS A DON'T CARE | AND, do not invert A, do not invert B 
	assign Dsel = 2'b01; //Enable ALU on data bus
	assign PCsel = 1'b1; //Pass A to PC
	assign SL = 1'b0;
	
	assign controlWord = {Psel, DA, SA, SB, Fsel, regW, ramW, Dsel, Bsel, PCsel, SL};
	
	assign nextState = 2'b00;
	
	assign K = {64'd0}; //THIS IS A DON'T CARE
	
endmodule
