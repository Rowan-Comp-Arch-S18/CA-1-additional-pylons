module ProgramCounter(PC, PC4, );