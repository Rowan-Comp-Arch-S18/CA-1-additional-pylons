module ROM_Pixel_Test(out, address);
   input[15:0] address;
   output reg[31:0] out;
   always @(address) begin
      case(address)
         16'd0: out = 32'b11010010100000000000000001010100; // MOVZ X20, 2
         16'd1: out = 32'b11010011011000001110001010010100; // LSL X20, X20, 56
         16'd2: out = 32'b10010001000000000000101010010101; // ADDI X21, X20, 2
         16'd3: out = 32'b10010001000010010111001010010110; // ADDI X22, X20, 604
         16'd4: out = 32'b11111000010000000000001010101010; // LDUR X10, [X21, 0]
         16'd5: out = 32'b10010010000000000000100101001010; // ANDI X10, X10, 2
         16'd6: out = 32'b10110100111111111111111110101010; // CBZ X10, -3
         16'd7: out = 32'b11111000010000000000001010101010; // LDUR X10, [X21, 0]
         16'd8: out = 32'b10010010000000000000010101001010; // ANDI X10, X10, 1
         16'd9: out = 32'b10110100111111111111111110101010; // CBZ X10, -3
         16'd10: out = 32'b11010010100110000000011000000000; // MOVZ X0, 49200
         16'd11: out = 32'b11010011011000001100000000000001; // LSL X1, X0, 48
         16'd12: out = 32'b11010010100000011001111000000000; // MOVZ X0, 3312
         16'd13: out = 32'b11010011011000001000000000000000; // LSL X0, X0, 32
         16'd14: out = 32'b10001011000000010000000000000001; // ADD X1, X0, X1
         16'd15: out = 32'b11010010100001111001100110000000; // MOVZ X0, 15564
         16'd16: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd17: out = 32'b10001011000000010000000000000001; // ADD X1, X0, X1
         16'd18: out = 32'b11010010100010101001111110000000; // MOVZ X0, 21756
         16'd19: out = 32'b10001011000000010000000000000001; // ADD X1, X0, X1
         16'd20: out = 32'b11111000000000000000001011000001; // STUR X1, [X22, 0]
         16'd21: out = 32'b10010001000000000000011011010110; // ADDI X22, X22, 1
         16'd22: out = 32'b11010001000100101101001011011001; // SUBI X25, X22, 1204
         16'd23: out = 32'b11001011000101000000001100111001; // SUB X25, X25, X20
         16'd24: out = 32'b10110101111111111111111101111001; // CBNZ X25, -5
         16'd25: out = 32'b11010010100000000000000010100101; // MOVZ X5, 5
         16'd26: out = 32'b11111000000000000000001010000101; // STUR X5, [X20, 0]
         16'd27: out = 32'b00010111111111111111111111111111; // B -1
         default: out = 32'b11010110000000000000001111100000; // BR XZR
      endcase
   end
endmodule
