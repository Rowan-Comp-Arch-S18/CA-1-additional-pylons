module ROM_Image_Display(out, address);
   input[15:0] address;
   output reg[31:0] out;
   always @(address) begin
      case(address)
         16'd0: out = 32'b11010010100000000000000001010100; // MOVZ X20, 2
         16'd1: out = 32'b11010011011000001110001010010100; // LSL X20, X20, 56
         16'd2: out = 32'b10010001000000000000101010010101; // ADDI X21, X20, 2
         16'd3: out = 32'b10010001000010010111001010010110; // ADDI X22, X20, 604
         16'd4: out = 32'b10001011000111110000001011000010; // ADD X2, X22, XZR
         16'd5: out = 32'b11111000010000000000001010100011; // LDUR X3, [X21, 0]
         16'd6: out = 32'b10010010000000000000100001100011; // ANDI X3, X3, 2
         16'd7: out = 32'b10110100111111111111111110100011; // CBZ X3, -3
         16'd8: out = 32'b11111000010000000000001010100011; // LDUR X3, [X21, 0]
         16'd9: out = 32'b10010010000000000000010001100011; // ANDI X3, X3, 1
         16'd10: out = 32'b10110100111111111111111110100011; // CBZ X3, -3
         16'd11: out = 32'b11010010100010100000101000000101; // MOVZ X5, 20560
         16'd12: out = 32'b10001011000010100000000010101010; // ADD X10, X5, X10
         16'd13: out = 32'b11010011011000000100000010100101; // LSL X5, X5, 16
         16'd14: out = 32'b10001011000010100000000010101010; // ADD X10, X5, X10
         16'd15: out = 32'b11010011011000000100000010100101; // LSL X5, X5, 16
         16'd16: out = 32'b10001011000010100000000010101010; // ADD X10, X5, X10
         16'd17: out = 32'b11010011011000000100000010100101; // LSL X5, X5, 16
         16'd18: out = 32'b10001011000010100000000010101010; // ADD X10, X5, X10
         16'd19: out = 32'b11010010100111001010001100000110; // MOVZ X6, 58648
         16'd20: out = 32'b10001011000010110000000011001011; // ADD X11, X6, X11
         16'd21: out = 32'b11010011011000000100000011000110; // LSL X6, X6, 16
         16'd22: out = 32'b10001011000010110000000011001011; // ADD X11, X6, X11
         16'd23: out = 32'b11010011011000000100000011000110; // LSL X6, X6, 16
         16'd24: out = 32'b10001011000010110000000011001011; // ADD X11, X6, X11
         16'd25: out = 32'b11010011011000000100000011000110; // LSL X6, X6, 16
         16'd26: out = 32'b10001011000010110000000011001011; // ADD X11, X6, X11
         16'd27: out = 32'b11010010100010101000101010000111; // MOVZ X7, 21588
         16'd28: out = 32'b10001011000011000000000011101100; // ADD X12, X7, X12
         16'd29: out = 32'b11010011011000000100000011100111; // LSL X7, X7, 16
         16'd30: out = 32'b10001011000011000000000011101100; // ADD X12, X7, X12
         16'd31: out = 32'b11010011011000000100000011100111; // LSL X7, X7, 16
         16'd32: out = 32'b10001011000011000000000011101100; // ADD X12, X7, X12
         16'd33: out = 32'b11010011011000000100000011100111; // LSL X7, X7, 16
         16'd34: out = 32'b10001011000011000000000011101100; // ADD X12, X7, X12
         16'd35: out = 32'b11010010100111110001111100001000; // MOVZ X8, 63736
         16'd36: out = 32'b10001011000011010000000100001101; // ADD X13, X8, X13
         16'd37: out = 32'b11010011011000000100000100001000; // LSL X8, X8, 16
         16'd38: out = 32'b10001011000011010000000100001101; // ADD X13, X8, X13
         16'd39: out = 32'b11010011011000000100000100001000; // LSL X8, X8, 16
         16'd40: out = 32'b10001011000011010000000100001101; // ADD X13, X8, X13
         16'd41: out = 32'b11010011011000000100000100001000; // LSL X8, X8, 16
         16'd42: out = 32'b10001011000011010000000100001101; // ADD X13, X8, X13
         16'd43: out = 32'b11010010100111111001111110001001; // MOVZ X9, 64764
         16'd44: out = 32'b10001011000011100000000100101110; // ADD X14, X9, X14
         16'd45: out = 32'b11010011011000000100000100101001; // LSL X9, X9, 16
         16'd46: out = 32'b10001011000011100000000100101110; // ADD X14, X9, X14
         16'd47: out = 32'b11010011011000000100000100101001; // LSL X9, X9, 16
         16'd48: out = 32'b10001011000011100000000100101110; // ADD X14, X9, X14
         16'd49: out = 32'b11010011011000000100000100101001; // LSL X9, X9, 16
         16'd50: out = 32'b10001011000011100000000100101110; // ADD X14, X9, X14
         16'd51: out = 32'b11010010100011001000110010001001; // MOVZ X9, 25700
         16'd52: out = 32'b10001011000011110000000100101111; // ADD X15, X9, X15
         16'd53: out = 32'b11010011011000000100000100101001; // LSL X9, X9, 16
         16'd54: out = 32'b10001011000011110000000100101111; // ADD X15, X9, X15
         16'd55: out = 32'b11010011011000000100000100101001; // LSL X9, X9, 16
         16'd56: out = 32'b10001011000011110000000100101111; // ADD X15, X9, X15
         16'd57: out = 32'b11010011011000000100000100101001; // LSL X9, X9, 16
         16'd58: out = 32'b10001011000011110000000100101111; // ADD X15, X9, X15
         16'd59: out = 32'b11010010100101001001010010001001; // MOVZ X9, 42148
         16'd60: out = 32'b10001011000100000000000100110000; // ADD X16, X9, X16
         16'd61: out = 32'b11010011011000000100000100101001; // LSL X9, X9, 16
         16'd62: out = 32'b10001011000100000000000100110000; // ADD X16, X9, X16
         16'd63: out = 32'b11010011011000000100000100101001; // LSL X9, X9, 16
         16'd64: out = 32'b10001011000100000000000100110000; // ADD X16, X9, X16
         16'd65: out = 32'b11010011011000000100000100101001; // LSL X9, X9, 16
         16'd66: out = 32'b10001011000100000000000100110000; // ADD X16, X9, X16
         16'd67: out = 32'b11010010100111010001110100001001; // MOVZ X9, 59624
         16'd68: out = 32'b10001011000100010000000100110001; // ADD X17, X9, X17
         16'd69: out = 32'b11010011011000000100000100101001; // LSL X9, X9, 16
         16'd70: out = 32'b10001011000100010000000100110001; // ADD X17, X9, X17
         16'd71: out = 32'b11010011011000000100000100101001; // LSL X9, X9, 16
         16'd72: out = 32'b10001011000100010000000100110001; // ADD X17, X9, X17
         16'd73: out = 32'b11010011011000000100000100101001; // LSL X9, X9, 16
         16'd74: out = 32'b10001011000100010000000100110001; // ADD X17, X9, X17
         16'd75: out = 32'b11010010100000001000000010001001; // MOVZ X9, 1028
         16'd76: out = 32'b10001011000100110000000100110011; // ADD X19, X9, X19
         16'd77: out = 32'b11010011011000000100000100101001; // LSL X9, X9, 16
         16'd78: out = 32'b10001011000100110000000100110011; // ADD X19, X9, X19
         16'd79: out = 32'b11010011011000000100000100101001; // LSL X9, X9, 16
         16'd80: out = 32'b10001011000100110000000100110011; // ADD X19, X9, X19
         16'd81: out = 32'b11010011011000000100000100101001; // LSL X9, X9, 16
         16'd82: out = 32'b10001011000100110000000100110011; // ADD X19, X9, X19
         16'd83: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd84: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd85: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd86: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd87: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd88: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd89: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd90: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd91: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd92: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd93: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd94: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd95: out = 32'b11110010100000000000000010000001; // MOVK X1, 4
         16'd96: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd97: out = 32'b11110010100010001000101010000001; // MOVK X1, 17492
         16'd98: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd99: out = 32'b10010001000000000001100001000010; // ADDI X2, X2, 6
         16'd100: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd101: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd102: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd103: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd104: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd105: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd106: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd107: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd108: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd109: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd110: out = 32'b11110010100010000000000000000001; // MOVK X1, 16384
         16'd111: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd112: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd113: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd114: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd115: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd116: out = 32'b10010001000000000001100001000010; // ADDI X2, X2, 6
         16'd117: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd118: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd119: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd120: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd121: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd122: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd123: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd124: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd125: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd126: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd127: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd128: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd129: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd130: out = 32'b11110010100000000000100000000001; // MOVK X1, 64
         16'd131: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd132: out = 32'b11110010100010000000101000000001; // MOVK X1, 16464
         16'd133: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd134: out = 32'b11110010100010100000101000000001; // MOVK X1, 20560
         16'd135: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd136: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd137: out = 32'b11010010100010000000101010000001; // MOVZ X1, 16468
         16'd138: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd139: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd140: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd141: out = 32'b11110010100000000000000010000001; // MOVK X1, 4
         16'd142: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd143: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd144: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd145: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd146: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd147: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd148: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd149: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd150: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd151: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd152: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd153: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd154: out = 32'b10010001000000000001100001000010; // ADDI X2, X2, 6
         16'd155: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd156: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd157: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd158: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd159: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd160: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd161: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd162: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd163: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd164: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd165: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd166: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd167: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd168: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd169: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd170: out = 32'b11110010100000000000101000000001; // MOVK X1, 80
         16'd171: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd172: out = 32'b11110010100100101001010010000001; // MOVK X1, 38052
         16'd173: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd174: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd175: out = 32'b11010010100010100000101010000001; // MOVZ X1, 20564
         16'd176: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd177: out = 32'b11110010100010000000000000000001; // MOVK X1, 16384
         16'd178: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd179: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd180: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd181: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd182: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd183: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd184: out = 32'b11111000000000000000000001010011; // STUR X19, [X2, 0]
         16'd185: out = 32'b10010001000000000001100001000010; // ADDI X2, X2, 6
         16'd186: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd187: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd188: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd189: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd190: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd191: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd192: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd193: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd194: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd195: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd196: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd197: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd198: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd199: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd200: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd201: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd202: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd203: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd204: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd205: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd206: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd207: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd208: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd209: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd210: out = 32'b11110010100010101001110100000001; // MOVK X1, 21736
         16'd211: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd212: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd213: out = 32'b11010010100111010001001010000001; // MOVZ X1, 59540
         16'd214: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd215: out = 32'b11110010100010100000000000000001; // MOVK X1, 20480
         16'd216: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd217: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd218: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd219: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd220: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd221: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd222: out = 32'b11111000000000000000000001010011; // STUR X19, [X2, 0]
         16'd223: out = 32'b10010001000000000001100001000010; // ADDI X2, X2, 6
         16'd224: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd225: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd226: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd227: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd228: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd229: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd230: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd231: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd232: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd233: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd234: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd235: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd236: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd237: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd238: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd239: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd240: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd241: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd242: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd243: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd244: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd245: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd246: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd247: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd248: out = 32'b11110010100000000000101000000001; // MOVK X1, 80
         16'd249: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd250: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd251: out = 32'b11010010100111010001010100000001; // MOVZ X1, 59560
         16'd252: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd253: out = 32'b11110010100010100000000000000001; // MOVK X1, 20480
         16'd254: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd255: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd256: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd257: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd258: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd259: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd260: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd261: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd262: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd263: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd264: out = 32'b11110010100000000000000010000001; // MOVK X1, 4
         16'd265: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd266: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd267: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd268: out = 32'b10010001000000000001100001000010; // ADDI X2, X2, 6
         16'd269: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd270: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd271: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd272: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd273: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd274: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd275: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd276: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd277: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd278: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd279: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd280: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd281: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd282: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd283: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd284: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd285: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd286: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd287: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd288: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd289: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd290: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd291: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd292: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd293: out = 32'b11110010100000000000100000000001; // MOVK X1, 64
         16'd294: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd295: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd296: out = 32'b11010010100101001001110100000001; // MOVZ X1, 42216
         16'd297: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd298: out = 32'b11110010100010101000000000000001; // MOVK X1, 21504
         16'd299: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd300: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd301: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd302: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd303: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd304: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd305: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd306: out = 32'b10010001000000000001100001000010; // ADDI X2, X2, 6
         16'd307: out = 32'b11010010100000010000000100000001; // MOVZ X1, 2056
         16'd308: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd309: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd310: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd311: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd312: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd313: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd314: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd315: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd316: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd317: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd318: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd319: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd320: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd321: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd322: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd323: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd324: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd325: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd326: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd327: out = 32'b11010010100010100001010010000001; // MOVZ X1, 20644
         16'd328: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd329: out = 32'b11110010100101001000101000000001; // MOVK X1, 42064
         16'd330: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd331: out = 32'b11110010100010000000000000000001; // MOVK X1, 16384
         16'd332: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd333: out = 32'b11110010100000000001010100000001; // MOVK X1, 168
         16'd334: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd335: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd336: out = 32'b10010001000000000001100001000010; // ADDI X2, X2, 6
         16'd337: out = 32'b11010010100000010000000100000001; // MOVZ X1, 2056
         16'd338: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd339: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd340: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd341: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd342: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd343: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd344: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd345: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd346: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd347: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd348: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd349: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd350: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd351: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd352: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd353: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd354: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd355: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd356: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd357: out = 32'b11010010100010000001001010000001; // MOVZ X1, 16532
         16'd358: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd359: out = 32'b11110010100101001001001010000001; // MOVK X1, 42132
         16'd360: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd361: out = 32'b11110010100100101000100000000001; // MOVK X1, 37952
         16'd362: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd363: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd364: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd365: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd366: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd367: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd368: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd369: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd370: out = 32'b11110010100000000000000010000001; // MOVK X1, 4
         16'd371: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd372: out = 32'b11110010100010101000101010000001; // MOVK X1, 21588
         16'd373: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd374: out = 32'b10010001000000000001100001000010; // ADDI X2, X2, 6
         16'd375: out = 32'b11010010100000010000000100000001; // MOVZ X1, 2056
         16'd376: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd377: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd378: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd379: out = 32'b11110010100000010000000010000001; // MOVK X1, 2052
         16'd380: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd381: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd382: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd383: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd384: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd385: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd386: out = 32'b11110010100000001000000100000001; // MOVK X1, 1032
         16'd387: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd388: out = 32'b11110010100010110000101100000001; // MOVK X1, 22616
         16'd389: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd390: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd391: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd392: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd393: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd394: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd395: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd396: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd397: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd398: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd399: out = 32'b11110010100000000000100000000001; // MOVK X1, 64
         16'd400: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd401: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd402: out = 32'b11010010100100101001110100000001; // MOVZ X1, 38120
         16'd403: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd404: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd405: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd406: out = 32'b11110010100111010000101010000001; // MOVK X1, 59476
         16'd407: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd408: out = 32'b11110010100000000000100000000001; // MOVK X1, 64
         16'd409: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd410: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd411: out = 32'b11010010100010000000000000000001; // MOVZ X1, 16384
         16'd412: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd413: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd414: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd415: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd416: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd417: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd418: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd419: out = 32'b10010001000000000001100001000010; // ADDI X2, X2, 6
         16'd420: out = 32'b11010010100000010000000100000001; // MOVZ X1, 2056
         16'd421: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd422: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd423: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd424: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd425: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd426: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd427: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd428: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd429: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd430: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd431: out = 32'b11110010100000010000001100000001; // MOVK X1, 2072
         16'd432: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd433: out = 32'b11110010100010110000101100000001; // MOVK X1, 22616
         16'd434: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd435: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd436: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd437: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd438: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd439: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd440: out = 32'b11110010100000000000100000000001; // MOVK X1, 64
         16'd441: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd442: out = 32'b11110010100010100001001010000001; // MOVK X1, 20628
         16'd443: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd444: out = 32'b11110010100111010001111100000001; // MOVK X1, 59640
         16'd445: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd446: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd447: out = 32'b11010010100111111001111110000001; // MOVZ X1, 64764
         16'd448: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd449: out = 32'b11110010100111110001111100000001; // MOVK X1, 63736
         16'd450: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd451: out = 32'b11110010100111010001001010000001; // MOVK X1, 59540
         16'd452: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd453: out = 32'b11110010100010100001001010000001; // MOVK X1, 20628
         16'd454: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd455: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd456: out = 32'b11010010100100101000000000000001; // MOVZ X1, 37888
         16'd457: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd458: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd459: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd460: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd461: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd462: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd463: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd464: out = 32'b10010001000000000001100001000010; // ADDI X2, X2, 6
         16'd465: out = 32'b11010010100000010000000100000001; // MOVZ X1, 2056
         16'd466: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd467: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd468: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd469: out = 32'b11110010100000010000101100000001; // MOVK X1, 2136
         16'd470: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd471: out = 32'b11110010100010110000101100000001; // MOVK X1, 22616
         16'd472: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd473: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd474: out = 32'b11010010100010110000000100000001; // MOVZ X1, 22536
         16'd475: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd476: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd477: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd478: out = 32'b11110010100000001000101010000001; // MOVK X1, 1108
         16'd479: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd480: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd481: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd482: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd483: out = 32'b11010010100000000000100000000001; // MOVZ X1, 64
         16'd484: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd485: out = 32'b11110010100010000000101000000001; // MOVK X1, 16464
         16'd486: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd487: out = 32'b11110010100010000000101000000001; // MOVK X1, 16464
         16'd488: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd489: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd490: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd491: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd492: out = 32'b11010010100111110001111100000001; // MOVZ X1, 63736
         16'd493: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd494: out = 32'b11110010100111110001110100000001; // MOVK X1, 63720
         16'd495: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd496: out = 32'b11110010100111010001001010000001; // MOVK X1, 59540
         16'd497: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd498: out = 32'b11110010100010101001001010000001; // MOVK X1, 21652
         16'd499: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd500: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd501: out = 32'b11010010100110101000101000000001; // MOVZ X1, 54352
         16'd502: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd503: out = 32'b11110010100000000000101000000001; // MOVK X1, 80
         16'd504: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd505: out = 32'b11110010100100100000100000000001; // MOVK X1, 36928
         16'd506: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd507: out = 32'b11110010100000000000101000000001; // MOVK X1, 80
         16'd508: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd509: out = 32'b10010001000000000001100001000010; // ADDI X2, X2, 6
         16'd510: out = 32'b11010010100000010000000100000001; // MOVZ X1, 2056
         16'd511: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd512: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd513: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd514: out = 32'b11110010100000000000000010000001; // MOVK X1, 4
         16'd515: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd516: out = 32'b11110010100000001000000100000001; // MOVK X1, 1032
         16'd517: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd518: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd519: out = 32'b11010010100000010000000010000001; // MOVZ X1, 2052
         16'd520: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd521: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd522: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd523: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd524: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd525: out = 32'b11110010100010000000000000000001; // MOVK X1, 16384
         16'd526: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd527: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd528: out = 32'b11010010100010000001001010000001; // MOVZ X1, 16532
         16'd529: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd530: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd531: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd532: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd533: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd534: out = 32'b11110010100010000001010010000001; // MOVK X1, 16548
         16'd535: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd536: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd537: out = 32'b11010010100111010001110010000001; // MOVZ X1, 59620
         16'd538: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd539: out = 32'b11110010100100101001110100000001; // MOVK X1, 38120
         16'd540: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd541: out = 32'b11110010100111010000101010000001; // MOVK X1, 59476
         16'd542: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd543: out = 32'b11110010100000000000101000000001; // MOVK X1, 80
         16'd544: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd545: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd546: out = 32'b11010010100111001001010010000001; // MOVZ X1, 58532
         16'd547: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd548: out = 32'b11110010100011001001010010000001; // MOVK X1, 25764
         16'd549: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd550: out = 32'b11110010100111001001010010000001; // MOVK X1, 58532
         16'd551: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd552: out = 32'b11110010100011001001010010000001; // MOVK X1, 25764
         16'd553: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd554: out = 32'b10010001000000000001100001000010; // ADDI X2, X2, 6
         16'd555: out = 32'b11010010100000010000000100000001; // MOVZ X1, 2056
         16'd556: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd557: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd558: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd559: out = 32'b11110010100000000000000010000001; // MOVK X1, 4
         16'd560: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd561: out = 32'b11110010100010101000101010000001; // MOVK X1, 21588
         16'd562: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd563: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd564: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd565: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd566: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd567: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd568: out = 32'b11110010100000001000100010000001; // MOVK X1, 1092
         16'd569: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd570: out = 32'b11110010100100101000100000000001; // MOVK X1, 37952
         16'd571: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd572: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd573: out = 32'b11010010100100100001001010000001; // MOVZ X1, 37012
         16'd574: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd575: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd576: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd577: out = 32'b11110010100101001001110100000001; // MOVK X1, 42216
         16'd578: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd579: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd580: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd581: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd582: out = 32'b11010010100111010000101000000001; // MOVZ X1, 59472
         16'd583: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd584: out = 32'b11110010100010000001001010000001; // MOVK X1, 16532
         16'd585: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd586: out = 32'b11110010100111010000100000000001; // MOVK X1, 59456
         16'd587: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd588: out = 32'b11110010100000000000110010000001; // MOVK X1, 100
         16'd589: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd590: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd591: out = 32'b11010010100101001001010010000001; // MOVZ X1, 42148
         16'd592: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd593: out = 32'b11110010100011001001010010000001; // MOVK X1, 25764
         16'd594: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd595: out = 32'b11110010100100100001010010000001; // MOVK X1, 37028
         16'd596: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd597: out = 32'b11110010100011001001010010000001; // MOVK X1, 25764
         16'd598: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd599: out = 32'b10010001000000000001100001000010; // ADDI X2, X2, 6
         16'd600: out = 32'b11010010100000010000000100000001; // MOVZ X1, 2056
         16'd601: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd602: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd603: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd604: out = 32'b11110010100000000000000010000001; // MOVK X1, 4
         16'd605: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd606: out = 32'b11110010100010101000000010000001; // MOVK X1, 21508
         16'd607: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd608: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd609: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd610: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd611: out = 32'b11110010100010001000101010000001; // MOVK X1, 17492
         16'd612: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd613: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd614: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd615: out = 32'b11110010100100101001001000000001; // MOVK X1, 38032
         16'd616: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd617: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd618: out = 32'b11010010100100101001001010000001; // MOVZ X1, 38036
         16'd619: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd620: out = 32'b11110010100100101001110100000001; // MOVK X1, 38120
         16'd621: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd622: out = 32'b11110010100111010001110010000001; // MOVK X1, 59620
         16'd623: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd624: out = 32'b11110010100100101001110100000001; // MOVK X1, 38120
         16'd625: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd626: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd627: out = 32'b11010010100111010001110100000001; // MOVZ X1, 59624
         16'd628: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd629: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd630: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd631: out = 32'b11110010100100101000000000000001; // MOVK X1, 37888
         16'd632: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd633: out = 32'b11110010100000000000110000000001; // MOVK X1, 96
         16'd634: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd635: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd636: out = 32'b11010010100101000000110010000001; // MOVZ X1, 41060
         16'd637: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd638: out = 32'b11110010100011001000110010000001; // MOVK X1, 25700
         16'd639: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd640: out = 32'b11110010100010100000110000000001; // MOVK X1, 20576
         16'd641: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd642: out = 32'b11110010100011001000110000000001; // MOVK X1, 25696
         16'd643: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd644: out = 32'b10010001000000000001100001000010; // ADDI X2, X2, 6
         16'd645: out = 32'b11010010100000010000000100000001; // MOVZ X1, 2056
         16'd646: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd647: out = 32'b11110010100000010000000010000001; // MOVK X1, 2052
         16'd648: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd649: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd650: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd651: out = 32'b11110010100010110000000010000001; // MOVK X1, 22532
         16'd652: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd653: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd654: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd655: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd656: out = 32'b11110010100010001000101010000001; // MOVK X1, 17492
         16'd657: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd658: out = 32'b11110010100000001000100010000001; // MOVK X1, 1092
         16'd659: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd660: out = 32'b11110010100100101001001000000001; // MOVK X1, 38032
         16'd661: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd662: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd663: out = 32'b11010010100100100001001000000001; // MOVZ X1, 37008
         16'd664: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd665: out = 32'b11110010100100101001110100000001; // MOVK X1, 38120
         16'd666: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd667: out = 32'b11110010100100101001101010000001; // MOVK X1, 38100
         16'd668: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd669: out = 32'b11110010100110101001110100000001; // MOVK X1, 54504
         16'd670: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd671: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd672: out = 32'b11010010100111010001110100000001; // MOVZ X1, 59624
         16'd673: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd674: out = 32'b11110010100111010001110010000001; // MOVK X1, 59620
         16'd675: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd676: out = 32'b11110010100010000000000000000001; // MOVK X1, 16384
         16'd677: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd678: out = 32'b11110010100000000000110010000001; // MOVK X1, 100
         16'd679: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd680: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd681: out = 32'b11010010100111000001010000000001; // MOVZ X1, 57504
         16'd682: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd683: out = 32'b11110010100011001001010000000001; // MOVK X1, 25760
         16'd684: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd685: out = 32'b11110010100111001000100000000001; // MOVK X1, 58432
         16'd686: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd687: out = 32'b11110010100011001001010010000001; // MOVK X1, 25764
         16'd688: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd689: out = 32'b10010001000000000001100001000010; // ADDI X2, X2, 6
         16'd690: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd691: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd692: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd693: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd694: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd695: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd696: out = 32'b11110010100010110000000010000001; // MOVK X1, 22532
         16'd697: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd698: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd699: out = 32'b11010010100000001000000000000001; // MOVZ X1, 1024
         16'd700: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd701: out = 32'b11110010100010101000101010000001; // MOVK X1, 21588
         16'd702: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd703: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd704: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd705: out = 32'b11110010100100101000101000000001; // MOVK X1, 37968
         16'd706: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd707: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd708: out = 32'b11010010100010100001001000000001; // MOVZ X1, 20624
         16'd709: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd710: out = 32'b11110010100100101001110010000001; // MOVK X1, 38116
         16'd711: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd712: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd713: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd714: out = 32'b11110010100100101001110100000001; // MOVK X1, 38120
         16'd715: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd716: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd717: out = 32'b11010010100111010001110100000001; // MOVZ X1, 59624
         16'd718: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd719: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd720: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd721: out = 32'b11110010100010101000000000000001; // MOVK X1, 21504
         16'd722: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd723: out = 32'b11110010100000000000110010000001; // MOVK X1, 100
         16'd724: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd725: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd726: out = 32'b11010010100101000001010000000001; // MOVZ X1, 41120
         16'd727: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd728: out = 32'b11110010100011001001010010000001; // MOVK X1, 25764
         16'd729: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd730: out = 32'b11110010100101000000101000000001; // MOVK X1, 41040
         16'd731: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd732: out = 32'b11110010100101001001110010000001; // MOVK X1, 42212
         16'd733: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd734: out = 32'b10010001000000000001100001000010; // ADDI X2, X2, 6
         16'd735: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd736: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd737: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd738: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd739: out = 32'b11110010100000000000000010000001; // MOVK X1, 4
         16'd740: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd741: out = 32'b11110010100010110000000010000001; // MOVK X1, 22532
         16'd742: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd743: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd744: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd745: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd746: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd747: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd748: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd749: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd750: out = 32'b11110010100000000000101000000001; // MOVK X1, 80
         16'd751: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd752: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd753: out = 32'b11010010100010000000100000000001; // MOVZ X1, 16448
         16'd754: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd755: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd756: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd757: out = 32'b11110010100010100000100000000001; // MOVK X1, 20544
         16'd758: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd759: out = 32'b11110010100010000001001010000001; // MOVK X1, 16532
         16'd760: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd761: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd762: out = 32'b11010010100101001001110010000001; // MOVZ X1, 42212
         16'd763: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd764: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd765: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd766: out = 32'b11110010100100101000000000000001; // MOVK X1, 37888
         16'd767: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd768: out = 32'b11110010100000100000101000000001; // MOVK X1, 4176
         16'd769: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd770: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd771: out = 32'b11010010100101001000110010000001; // MOVZ X1, 42084
         16'd772: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd773: out = 32'b11110010100011000000110010000001; // MOVK X1, 24676
         16'd774: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd775: out = 32'b11110010100011000000000000000001; // MOVK X1, 24576
         16'd776: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd777: out = 32'b11110010100101001001001010000001; // MOVK X1, 42132
         16'd778: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd779: out = 32'b10010001000000000001100001000010; // ADDI X2, X2, 6
         16'd780: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd781: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd782: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd783: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd784: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd785: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd786: out = 32'b11110010100010101000100010000001; // MOVK X1, 21572
         16'd787: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd788: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd789: out = 32'b11010010100010110000101100000001; // MOVZ X1, 22616
         16'd790: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd791: out = 32'b11110010100010110000000010000001; // MOVK X1, 22532
         16'd792: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd793: out = 32'b11110010100000000000101010000001; // MOVK X1, 84
         16'd794: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd795: out = 32'b11110010100000000000101000000001; // MOVK X1, 80
         16'd796: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd797: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd798: out = 32'b11010010100010000000100000000001; // MOVZ X1, 16448
         16'd799: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd800: out = 32'b11110010100100101000100000000001; // MOVK X1, 37952
         16'd801: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd802: out = 32'b11110010100010000001001010000001; // MOVK X1, 16532
         16'd803: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd804: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd805: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd806: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd807: out = 32'b11010010100111010001110010000001; // MOVZ X1, 59620
         16'd808: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd809: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd810: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd811: out = 32'b11110010100100101001001000000001; // MOVK X1, 38032
         16'd812: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd813: out = 32'b11110010100010101001010100000001; // MOVK X1, 21672
         16'd814: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd815: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd816: out = 32'b11010010100101001001001000000001; // MOVZ X1, 42128
         16'd817: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd818: out = 32'b11110010100000000000101000000001; // MOVK X1, 80
         16'd819: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd820: out = 32'b11110010100100100000101000000001; // MOVK X1, 36944
         16'd821: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd822: out = 32'b11110010100010101001001010000001; // MOVK X1, 21652
         16'd823: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd824: out = 32'b10010001000000000001100001000010; // ADDI X2, X2, 6
         16'd825: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd826: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd827: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd828: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd829: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd830: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd831: out = 32'b11110010100000001000101010000001; // MOVK X1, 1108
         16'd832: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd833: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd834: out = 32'b11010010100010110000101100000001; // MOVZ X1, 22616
         16'd835: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd836: out = 32'b11110010100010110000000010000001; // MOVK X1, 22532
         16'd837: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd838: out = 32'b11110010100000000000101010000001; // MOVK X1, 84
         16'd839: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd840: out = 32'b11110010100000000000101000000001; // MOVK X1, 80
         16'd841: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd842: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd843: out = 32'b11010010100010000000100000000001; // MOVZ X1, 16448
         16'd844: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd845: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd846: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd847: out = 32'b11110010100100101001010010000001; // MOVK X1, 38052
         16'd848: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd849: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd850: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd851: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd852: out = 32'b11010010100100101001110010000001; // MOVZ X1, 38116
         16'd853: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd854: out = 32'b11110010100111001001110100000001; // MOVK X1, 58600
         16'd855: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd856: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd857: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd858: out = 32'b11110010100010100000101010000001; // MOVK X1, 20564
         16'd859: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd860: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd861: out = 32'b11010010100111001001001010000001; // MOVZ X1, 58516
         16'd862: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd863: out = 32'b11110010100010100000100000000001; // MOVK X1, 20544
         16'd864: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd865: out = 32'b11110010100111001001001010000001; // MOVK X1, 58516
         16'd866: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd867: out = 32'b11110010100010101001110010000001; // MOVK X1, 21732
         16'd868: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd869: out = 32'b10010001000000000001100001000010; // ADDI X2, X2, 6
         16'd870: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd871: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd872: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd873: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd874: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd875: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd876: out = 32'b11110010100000000000000010000001; // MOVK X1, 4
         16'd877: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd878: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd879: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd880: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd881: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd882: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd883: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd884: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd885: out = 32'b11110010100000000000101000000001; // MOVK X1, 80
         16'd886: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd887: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd888: out = 32'b11010010100010000000100000000001; // MOVZ X1, 16448
         16'd889: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd890: out = 32'b11110010100100101001001000000001; // MOVK X1, 38032
         16'd891: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd892: out = 32'b11110010100100101001110100000001; // MOVK X1, 38120
         16'd893: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd894: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd895: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd896: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd897: out = 32'b11010010100111010001110100000001; // MOVZ X1, 59624
         16'd898: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd899: out = 32'b11110010100101001000100000000001; // MOVK X1, 42048
         16'd900: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd901: out = 32'b11110010100010100000101000000001; // MOVK X1, 20560
         16'd902: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd903: out = 32'b11110010100000100000001000000001; // MOVK X1, 4112
         16'd904: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd905: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd906: out = 32'b11010010100010100000101000000001; // MOVZ X1, 20560
         16'd907: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd908: out = 32'b11110010100000100000101010000001; // MOVK X1, 4180
         16'd909: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd910: out = 32'b11110010100101010001010010000001; // MOVK X1, 43172
         16'd911: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd912: out = 32'b11110010100101001001010010000001; // MOVK X1, 42148
         16'd913: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd914: out = 32'b10010001000000000001100001000010; // ADDI X2, X2, 6
         16'd915: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd916: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd917: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd918: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd919: out = 32'b11110010100010110000101100000001; // MOVK X1, 22616
         16'd920: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd921: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd922: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd923: out = 32'b11110010100000000000101000000001; // MOVK X1, 80
         16'd924: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd925: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd926: out = 32'b11010010100010000000100000000001; // MOVZ X1, 16448
         16'd927: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd928: out = 32'b11110010100100100001001010000001; // MOVK X1, 37012
         16'd929: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd930: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd931: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd932: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd933: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd934: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd935: out = 32'b11010010100111010001010010000001; // MOVZ X1, 59556
         16'd936: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd937: out = 32'b11110010100100101000000000000001; // MOVK X1, 37888
         16'd938: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd939: out = 32'b11110010100010100000101000000001; // MOVK X1, 20560
         16'd940: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd941: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd942: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd943: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd944: out = 32'b11010010100010100000101000000001; // MOVZ X1, 20560
         16'd945: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd946: out = 32'b11110010100000100000101000000001; // MOVK X1, 4176
         16'd947: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd948: out = 32'b11110010100010101000101010000001; // MOVK X1, 21588
         16'd949: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd950: out = 32'b11110010100101001001010010000001; // MOVK X1, 42148
         16'd951: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd952: out = 32'b10010001000000000001100001000010; // ADDI X2, X2, 6
         16'd953: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd954: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd955: out = 32'b11010010100000001000000000000001; // MOVZ X1, 1024
         16'd956: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd957: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd958: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd959: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd960: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd961: out = 32'b11110010100000000000100000000001; // MOVK X1, 64
         16'd962: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd963: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd964: out = 32'b11010010100010000000000000000001; // MOVZ X1, 16384
         16'd965: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd966: out = 32'b11110010100010000001001010000001; // MOVK X1, 16532
         16'd967: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd968: out = 32'b11110010100111001001110100000001; // MOVK X1, 58600
         16'd969: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd970: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd971: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd972: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd973: out = 32'b11010010100101001001010100000001; // MOVZ X1, 42152
         16'd974: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd975: out = 32'b11110010100111111001111110000001; // MOVK X1, 64764
         16'd976: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd977: out = 32'b11110010100111111001111110000001; // MOVK X1, 64764
         16'd978: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd979: out = 32'b11110010100111111001111110000001; // MOVK X1, 64764
         16'd980: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd981: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd982: out = 32'b11010010100111111001111110000001; // MOVZ X1, 64764
         16'd983: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd984: out = 32'b11110010100101110001110100000001; // MOVK X1, 47336
         16'd985: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd986: out = 32'b11110010100111010001010100000001; // MOVK X1, 59560
         16'd987: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd988: out = 32'b11110010100101010001111100000001; // MOVK X1, 43256
         16'd989: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd990: out = 32'b10010001000000000001100001000010; // ADDI X2, X2, 6
         16'd991: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd992: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd993: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd994: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd995: out = 32'b11010010100010000000000000000001; // MOVZ X1, 16384
         16'd996: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd997: out = 32'b11110010100000000000100000000001; // MOVK X1, 64
         16'd998: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd999: out = 32'b11110010100100101001110010000001; // MOVK X1, 38116
         16'd1000: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1001: out = 32'b11110010100111010001010010000001; // MOVK X1, 59556
         16'd1002: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1003: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1004: out = 32'b11010010100010100000101010000001; // MOVZ X1, 20564
         16'd1005: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1006: out = 32'b11110010100010101000101100000001; // MOVK X1, 21592
         16'd1007: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1008: out = 32'b11110010100011010000110100000001; // MOVK X1, 26728
         16'd1009: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1010: out = 32'b11110010100011010001010100000001; // MOVK X1, 26792
         16'd1011: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1012: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1013: out = 32'b11010010100101011001010110000001; // MOVZ X1, 44204
         16'd1014: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1015: out = 32'b11110010100101111001011110000001; // MOVK X1, 48316
         16'd1016: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1017: out = 32'b11110010100111111001111110000001; // MOVK X1, 64764
         16'd1018: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1019: out = 32'b11110010100111111001111110000001; // MOVK X1, 64764
         16'd1020: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1021: out = 32'b10010001000000000001100001000010; // ADDI X2, X2, 6
         16'd1022: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1023: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1024: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1025: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1026: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd1027: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1028: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1029: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1030: out = 32'b11110010100000000000100000000001; // MOVK X1, 64
         16'd1031: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1032: out = 32'b11110010100010000001001010000001; // MOVK X1, 16532
         16'd1033: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1034: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1035: out = 32'b11010010100010101000000000000001; // MOVZ X1, 21504
         16'd1036: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1037: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1038: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1039: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1040: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1041: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1042: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1043: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1044: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd1045: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1046: out = 32'b11110010100000000000000010000001; // MOVK X1, 4
         16'd1047: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1048: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1049: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1050: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1051: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1052: out = 32'b10010001000000000001100001000010; // ADDI X2, X2, 6
         16'd1053: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1054: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1055: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1056: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1057: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd1058: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1059: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1060: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1061: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1062: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1063: out = 32'b11110010100010100001010010000001; // MOVK X1, 20644
         16'd1064: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1065: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1066: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1067: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1068: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1069: out = 32'b10010001000000000001100001000010; // ADDI X2, X2, 6
         16'd1070: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1071: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1072: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1073: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1074: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd1075: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1076: out = 32'b11110010100000000000100000000001; // MOVK X1, 64
         16'd1077: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1078: out = 32'b11110010100010100001001010000001; // MOVK X1, 20628
         16'd1079: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1080: out = 32'b11110010100101001001010010000001; // MOVK X1, 42148
         16'd1081: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1082: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1083: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1084: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1085: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1086: out = 32'b10010001000000000001100001000010; // ADDI X2, X2, 6
         16'd1087: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1088: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1089: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1090: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1091: out = 32'b11010010100000000000101000000001; // MOVZ X1, 80
         16'd1092: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1093: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd1094: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1095: out = 32'b11110010100100101001010010000001; // MOVK X1, 38052
         16'd1096: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1097: out = 32'b11110010100111001001001010000001; // MOVK X1, 58516
         16'd1098: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1099: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1100: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1101: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1102: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1103: out = 32'b10010001000000000001100001000010; // ADDI X2, X2, 6
         16'd1104: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1105: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1106: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1107: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1108: out = 32'b11010010100101001001110100000001; // MOVZ X1, 42216
         16'd1109: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1110: out = 32'b11110010100111010001010010000001; // MOVK X1, 59556
         16'd1111: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1112: out = 32'b11110010100100101001010010000001; // MOVK X1, 38052
         16'd1113: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1114: out = 32'b11110010100111010000101000000001; // MOVK X1, 59472
         16'd1115: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1116: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1117: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1118: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1119: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1120: out = 32'b10010001000000000001100001000010; // ADDI X2, X2, 6
         16'd1121: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1122: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1123: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1124: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1125: out = 32'b11010010100000000001110100000001; // MOVZ X1, 232
         16'd1126: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1127: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd1128: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1129: out = 32'b11110010100101001001110100000001; // MOVK X1, 42216
         16'd1130: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1131: out = 32'b11110010100101010000000000000001; // MOVK X1, 43008
         16'd1132: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1133: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1134: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1135: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1136: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1137: out = 32'b10010001000000000001100001000010; // ADDI X2, X2, 6
         16'd1138: out = 32'b11010010100000000000000010100101; // MOVZ X5, 5
         16'd1139: out = 32'b11111000000000000000001010000101; // STUR X5, [X20, 0]
         16'd1140: out = 32'b00010111111111111111111111111111; // B -1
         default: out = 32'b11010110000000000000001111100000; // BR XZR
      endcase
   end
endmodule
