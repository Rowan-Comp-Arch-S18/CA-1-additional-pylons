module ROM_Flippy_Bit(out, address);
   input[15:0] address;
   output reg[31:0] out;
   always @(address) begin
      case(address)
         // InitAddresses: // ***** Create the address locations in ram - start at 8
         16'd0: out = 32'b11010010100000000010000000000001; // MOVZ X1, 256 // Blank RAM
         // IA-ClearRAM:
         16'd1: out = 32'b11010001000000000000010000100010; // SUBI X2, X1, 1
         16'd2: out = 32'b11111000000000000000000001011111; // STUR XZR, [X2, 0]
         16'd3: out = 32'b11010001000000000000010000100001; // SUBI X1, X1, 1
         16'd4: out = 32'b10110101111111111111111110000001; // CBNZ X1, IA-ClearRAM
         16'd5: out = 32'b11010010100000000000000001000000; // MOVZ X0, 2 // GPU
         16'd6: out = 32'b11010011011000001110000000000000; // LSL X0, X0, 56 // Control - 8
         16'd7: out = 32'b11111000000000001000001111100000; // STUR X0, [XZR, 8]
         16'd8: out = 32'b10010001000000000000100000000000; // ADDI X0, X0, 2 // Status - 9
         16'd9: out = 32'b11111000000000001001001111100000; // STUR X0, [XZR, 9]
         16'd10: out = 32'b10010001000010010110100000000000; // ADDI X0, X0, 602 // Top of screen - 10 - 480 locations
         16'd11: out = 32'b11111000000000001010001111100000; // STUR X0, [XZR, 10]
         16'd12: out = 32'b10010001000001111000000000000000; // ADDI X0, X0, 480 // Dark blue sky - 11 - 50 locations
         16'd13: out = 32'b11111000000000001011001111100000; // STUR X0, [XZR, 11]
         16'd14: out = 32'b10010001000000001100100000000000; // ADDI X0, X0, 50 // Ground - 12 - 70 locations
         16'd15: out = 32'b11111000000000001100001111100000; // STUR X0, [XZR, 12] // End of GPU addresses
         16'd16: out = 32'b11010010100000000000010000000001; // MOVZ X1, 32 // Counter
         // InitAlienData:
         16'd17: out = 32'b11111000000010111111000000111111; // STUR XZR, [X1, 191] // Start of Aliens - starts at 192 actually, just offset by the counter starting at 32
         16'd18: out = 32'b11010001000000000000010000100001; // SUBI X1, X1, 1
         16'd19: out = 32'b10110101111111111111111110100001; // CBNZ X1, InitAlienData // 32 Alien data 63=valid, 23-16=x, 15-8=y, 7-0=code
         16'd20: out = 32'b11111000000011111010001111111111; // STUR XZR, [XZR, 250] // Current score
         16'd21: out = 32'b11111000000011111011001111111111; // STUR XZR, [XZR, 251] // High score
         16'd22: out = 32'b11111000000011111100001111111111; // STUR XZR, [XZR, 252] // The current input
         16'd23: out = 32'b11111000000011111101001111111111; // STUR XZR, [XZR, 253] // The last input
         16'd24: out = 32'b11010010100000000000000000100000; // MOVZ X0, 1 // Keyboard
         16'd25: out = 32'b11010011011000001110000000000000; // LSL X0, X0, 56 // First keyboard register - 254
         16'd26: out = 32'b11111000000011111110001111100000; // STUR X0, [XZR, 254]
         16'd27: out = 32'b11010010100000000000000000100000; // MOVZ X0, 1 // Alien 1
         16'd28: out = 32'b11010011011000001011110000000000; // LSL X0, X0, 47
         16'd29: out = 32'b11110010100000000000000000000000; // MOVK X0, 0
         16'd30: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd31: out = 32'b11110010100001011010111010100000; // MOVK X0, 11637
         16'd32: out = 32'b11111000000011001000001111100000; // STUR X0, [XZR, 200]
         16'd33: out = 32'b11010010100000000000000000100000; // MOVZ X0, 1 // Alien 2
         16'd34: out = 32'b11010011011000001011110000000000; // LSL X0, X0, 47
         16'd35: out = 32'b11110010100000000000000010100000; // MOVK X0, 5
         16'd36: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd37: out = 32'b11110010100000101001101100000000; // MOVK X0, 5336
         16'd38: out = 32'b11111000000011001001001111100000; // STUR X0, [XZR, 201]
         16'd39: out = 32'b11010010100000000000000000100000; // MOVZ X0, 1 // Alien 3
         16'd40: out = 32'b11010011011000001011110000000000; // LSL X0, X0, 47
         16'd41: out = 32'b11110010100000000000000011100000; // MOVK X0, 7
         16'd42: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd43: out = 32'b11110010100001000000010101000000; // MOVK X0, 8234
         16'd44: out = 32'b11111000000011001010001111100000; // STUR X0, [XZR, 202]
         16'd45: out = 32'b00010100000000000000000000000000; // B InitColors // Next initialization step
         //
         // InitColors: // ***** Create the colors in ram - start at 0
         16'd46: out = 32'b11010010100111111001111110000000; // MOVZ X0, 64764 // White - 0
         16'd47: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd48: out = 32'b11110010100111111001111110000000; // MOVK X0, 64764
         16'd49: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd50: out = 32'b11110010100111111001111110000000; // MOVK X0, 64764
         16'd51: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd52: out = 32'b11110010100111111001111110000000; // MOVK X0, 64764
         16'd53: out = 32'b11111000000000000000001111100000; // STUR X0, [XZR, 0]
         16'd54: out = 32'b11010010100101011001010110000000; // MOVZ X0, 44204 // Light Blue - 1
         16'd55: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd56: out = 32'b11110010100101011001010110000000; // MOVK X0, 44204
         16'd57: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd58: out = 32'b11110010100101011001010110000000; // MOVK X0, 44204
         16'd59: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd60: out = 32'b11110010100101011001010110000000; // MOVK X0, 44204
         16'd61: out = 32'b11111000000000000001001111100000; // STUR X0, [XZR, 1]
         16'd62: out = 32'b11010010100101011001010110000000; // MOVZ X0, 44204 // Dark Blue - 2 - override to light blue
         16'd63: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd64: out = 32'b11110010100101011001010110000000; // MOVK X0, 44204
         16'd65: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd66: out = 32'b11110010100101011001010110000000; // MOVK X0, 44204
         16'd67: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd68: out = 32'b11110010100101011001010110000000; // MOVK X0, 44204
         16'd69: out = 32'b11111000000000000010001111100000; // STUR X0, [XZR, 2]
         16'd70: out = 32'b11010010100100100001001000000000; // MOVZ X0, 37008 // Brown - 3
         16'd71: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd72: out = 32'b11110010100100100001001000000000; // MOVK X0, 37008
         16'd73: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd74: out = 32'b11110010100100100001001000000000; // MOVK X0, 37008
         16'd75: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd76: out = 32'b11110010100100100001001000000000; // MOVK X0, 37008
         16'd77: out = 32'b11111000000000000011001111100000; // STUR X0, [XZR, 3]
         16'd78: out = 32'b11010010100111100001111000000000; // MOVZ X0, 61680 // Yellow - 4
         16'd79: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd80: out = 32'b11110010100111100001111000000000; // MOVK X0, 61680
         16'd81: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd82: out = 32'b11110010100111100001111000000000; // MOVK X0, 61680
         16'd83: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd84: out = 32'b11110010100111100001111000000000; // MOVK X0, 61680
         16'd85: out = 32'b11111000000000000100001111100000; // STUR X0, [XZR, 4]
         16'd86: out = 32'b11010010100110000001100000000000; // MOVZ X0, 49344 // Red - 5
         16'd87: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd88: out = 32'b11110010100110000001100000000000; // MOVK X0, 49344
         16'd89: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd90: out = 32'b11110010100110000001100000000000; // MOVK X0, 49344
         16'd91: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd92: out = 32'b11110010100110000001100000000000; // MOVK X0, 49344
         16'd93: out = 32'b11111000000000000101001111100000; // STUR X0, [XZR, 5]
         16'd94: out = 32'b00010100000000000000000000000000; // B InitBitmasks // Next initialization step
         //
         // InitBitmasks: // ***** Create the bitmasks for the text in ram - start at 16 - access with index << 3 + 16
         16'd95: out = 32'b11010010100111111000000000000000; // MOVZ X0, 64512 // Character 0
         16'd96: out = 32'b11111000000000010000001111100000; // STUR X0, [XZR, 16]
         16'd97: out = 32'b11010010100000000001111110000000; // MOVZ X0, 252
         16'd98: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd99: out = 32'b11110010100000000001111110000000; // MOVK X0, 252
         16'd100: out = 32'b11111000000000010001001111100000; // STUR X0, [XZR, 17]
         16'd101: out = 32'b11111000000000010010001111100000; // STUR X0, [XZR, 18]
         16'd102: out = 32'b11111000000000010011001111100000; // STUR X0, [XZR, 19]
         16'd103: out = 32'b11010010100111111000000000000000; // MOVZ X0, 64512
         16'd104: out = 32'b11111000000000010100001111100000; // STUR X0, [XZR, 20]
         16'd105: out = 32'b11010010100111111000000000000000; // MOVZ X0, 64512 // Character 1
         16'd106: out = 32'b11111000000000011000001111100000; // STUR X0, [XZR, 24]
         16'd107: out = 32'b11111000000000011001001111100000; // STUR X0, [XZR, 25]
         16'd108: out = 32'b11111000000000011010001111100000; // STUR X0, [XZR, 26]
         16'd109: out = 32'b11111000000000011011001111100000; // STUR X0, [XZR, 27]
         16'd110: out = 32'b11111000000000011100001111100000; // STUR X0, [XZR, 28]
         16'd111: out = 32'b11010010100000000001111110000000; // MOVZ X0, 252 // Character 2
         16'd112: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd113: out = 32'b11110010100111111000000000000000; // MOVK X0, 64512
         16'd114: out = 32'b11111000000000100000001111100000; // STUR X0, [XZR, 32]
         16'd115: out = 32'b11010010100000000001111110000000; // MOVZ X0, 252
         16'd116: out = 32'b11111000000000100001001111100000; // STUR X0, [XZR, 33]
         16'd117: out = 32'b11010010100111111000000000000000; // MOVZ X0, 64512
         16'd118: out = 32'b11111000000000100010001111100000; // STUR X0, [XZR, 34]
         16'd119: out = 32'b11010010100000000001111110000000; // MOVZ X0, 252
         16'd120: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd121: out = 32'b11111000000000100011001111100000; // STUR X0, [XZR, 35]
         16'd122: out = 32'b11110010100111111001111110000000; // MOVK X0, 64764
         16'd123: out = 32'b11111000000000100100001111100000; // STUR X0, [XZR, 36]
         16'd124: out = 32'b11010010100000000001111110000000; // MOVZ X0, 252 // Character 3
         16'd125: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd126: out = 32'b11110010100111111000000000000000; // MOVK X0, 64512
         16'd127: out = 32'b11111000000000101000001111100000; // STUR X0, [XZR, 40]
         16'd128: out = 32'b11111000000000101010001111100000; // STUR X0, [XZR, 42]
         16'd129: out = 32'b11111000000000101100001111100000; // STUR X0, [XZR, 44]
         16'd130: out = 32'b11010010100000000001111110000000; // MOVZ X0, 252
         16'd131: out = 32'b11111000000000101001001111100000; // STUR X0, [XZR, 41]
         16'd132: out = 32'b11111000000000101011001111100000; // STUR X0, [XZR, 43]
         16'd133: out = 32'b11010010100000000001111110000000; // MOVZ X0, 252 // Character 4
         16'd134: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd135: out = 32'b11110010100000000001111110000000; // MOVK X0, 252
         16'd136: out = 32'b11111000000000110000001111100000; // STUR X0, [XZR, 48]
         16'd137: out = 32'b11111000000000110001001111100000; // STUR X0, [XZR, 49]
         16'd138: out = 32'b11110010100111111001111110000000; // MOVK X0, 64764
         16'd139: out = 32'b11111000000000110010001111100000; // STUR X0, [XZR, 50]
         16'd140: out = 32'b11010010100000000001111110000000; // MOVZ X0, 252
         16'd141: out = 32'b11111000000000110011001111100000; // STUR X0, [XZR, 51]
         16'd142: out = 32'b11111000000000110100001111100000; // STUR X0, [XZR, 52]
         16'd143: out = 32'b11010010100000000001111110000000; // MOVZ X0, 252 // Character 5
         16'd144: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd145: out = 32'b11110010100111111001111110000000; // MOVK X0, 64764
         16'd146: out = 32'b11111000000000111000001111100000; // STUR X0, [XZR, 56]
         16'd147: out = 32'b11010010100000000001111110000000; // MOVZ X0, 252
         16'd148: out = 32'b11111000000000111011001111100000; // STUR X0, [XZR, 59]
         16'd149: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd150: out = 32'b11110010100000000000000000000000; // MOVK X0, 0
         16'd151: out = 32'b11111000000000111001001111100000; // STUR X0, [XZR, 57]
         16'd152: out = 32'b11010010100000000001111110000000; // MOVZ X0, 252
         16'd153: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd154: out = 32'b11110010100111111000000000000000; // MOVK X0, 64512
         16'd155: out = 32'b11111000000000111010001111100000; // STUR X0, [XZR, 58]
         16'd156: out = 32'b11111000000000111100001111100000; // STUR X0, [XZR, 60]
         16'd157: out = 32'b11010010100111111001111110000000; // MOVZ X0, 64764 // Character 6
         16'd158: out = 32'b11111000000001000000001111100000; // STUR X0, [XZR, 64]
         16'd159: out = 32'b11010011011000000010000000000000; // LSL X0, X0, 8
         16'd160: out = 32'b11111000000001000010001111100000; // STUR X0, [XZR, 66]
         16'd161: out = 32'b11010010100000000001111110000000; // MOVZ X0, 252
         16'd162: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd163: out = 32'b11111000000001000001001111100000; // STUR X0, [XZR, 65]
         16'd164: out = 32'b11110010100000000001111110000000; // MOVK X0, 252
         16'd165: out = 32'b11111000000001000011001111100000; // STUR X0, [XZR, 67]
         16'd166: out = 32'b11010010100111111000000000000000; // MOVZ X0, 64512
         16'd167: out = 32'b11111000000001000100001111100000; // STUR X0, [XZR, 68]
         16'd168: out = 32'b11010010100000000001111110000000; // MOVZ X0, 252 // Character 7
         16'd169: out = 32'b11111000000001001001001111100000; // STUR X0, [XZR, 73]
         16'd170: out = 32'b11010011011000000010000000000000; // LSL X0, X0, 8
         16'd171: out = 32'b11111000000001001010001111100000; // STUR X0, [XZR, 74]
         16'd172: out = 32'b11111000000001001011001111100000; // STUR X0, [XZR, 75]
         16'd173: out = 32'b11010011011000000010000000000000; // LSL X0, X0, 8
         16'd174: out = 32'b11111000000001001100001111100000; // STUR X0, [XZR, 76]
         16'd175: out = 32'b11110010100111111001111110000000; // MOVK X0, 64764
         16'd176: out = 32'b11111000000001001000001111100000; // STUR X0, [XZR, 72]
         16'd177: out = 32'b11010010100111111000000000000000; // MOVZ X0, 64512 // Character 8
         16'd178: out = 32'b11111000000001010000001111100000; // STUR X0, [XZR, 80]
         16'd179: out = 32'b11111000000001010010001111100000; // STUR X0, [XZR, 82]
         16'd180: out = 32'b11111000000001010100001111100000; // STUR X0, [XZR, 84]
         16'd181: out = 32'b11010010100000000001111110000000; // MOVZ X0, 252
         16'd182: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd183: out = 32'b11110010100000000001111110000000; // MOVK X0, 252
         16'd184: out = 32'b11111000000001010001001111100000; // STUR X0, [XZR, 81]
         16'd185: out = 32'b11111000000001010011001111100000; // STUR X0, [XZR, 83]
         16'd186: out = 32'b11010010100111111000000000000000; // MOVZ X0, 64512 // Character 9
         16'd187: out = 32'b11111000000001011000001111100000; // STUR X0, [XZR, 88]
         16'd188: out = 32'b11010010100000000001111110000000; // MOVZ X0, 252
         16'd189: out = 32'b11111000000001011011001111100000; // STUR X0, [XZR, 91]
         16'd190: out = 32'b11111000000001011100001111100000; // STUR X0, [XZR, 92]
         16'd191: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd192: out = 32'b11110010100000000001111110000000; // MOVK X0, 252
         16'd193: out = 32'b11111000000001011001001111100000; // STUR X0, [XZR, 89]
         16'd194: out = 32'b11010010100111111001111110000000; // MOVZ X0, 64764
         16'd195: out = 32'b11111000000001011010001111100000; // STUR X0, [XZR, 90]
         16'd196: out = 32'b11010010100111111000000000000000; // MOVZ X0, 64512 // Character A
         16'd197: out = 32'b11111000000001100000001111100000; // STUR X0, [XZR, 96]
         16'd198: out = 32'b11111000000001100001001111100000; // STUR X0, [XZR, 97]
         16'd199: out = 32'b11010010100000000001111110000000; // MOVZ X0, 252
         16'd200: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd201: out = 32'b11110010100000000001111110000000; // MOVK X0, 252
         16'd202: out = 32'b11111000000001100010001111100000; // STUR X0, [XZR, 98]
         16'd203: out = 32'b11111000000001100100001111100000; // STUR X0, [XZR, 100]
         16'd204: out = 32'b11110010100111111001111110000000; // MOVK X0, 64764
         16'd205: out = 32'b11111000000001100011001111100000; // STUR X0, [XZR, 99]
         16'd206: out = 32'b11010010100000000001111110000000; // MOVZ X0, 252 // Character B
         16'd207: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd208: out = 32'b11110010100111111000000000000000; // MOVK X0, 64512
         16'd209: out = 32'b11111000000001101000001111100000; // STUR X0, [XZR, 104]
         16'd210: out = 32'b11111000000001101010001111100000; // STUR X0, [XZR, 106]
         16'd211: out = 32'b11111000000001101100001111100000; // STUR X0, [XZR, 108]
         16'd212: out = 32'b11110010100000000001111110000000; // MOVK X0, 252
         16'd213: out = 32'b11111000000001101001001111100000; // STUR X0, [XZR, 105]
         16'd214: out = 32'b11111000000001101011001111100000; // STUR X0, [XZR, 107]
         16'd215: out = 32'b11010010100111111001111110000000; // MOVZ X0, 64764 // Character C
         16'd216: out = 32'b11111000000001110000001111100000; // STUR X0, [XZR, 112]
         16'd217: out = 32'b11111000000001110100001111100000; // STUR X0, [XZR, 116]
         16'd218: out = 32'b11010010100000000001111110000000; // MOVZ X0, 252
         16'd219: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd220: out = 32'b11111000000001110001001111100000; // STUR X0, [XZR, 113]
         16'd221: out = 32'b11111000000001110010001111100000; // STUR X0, [XZR, 114]
         16'd222: out = 32'b11111000000001110011001111100000; // STUR X0, [XZR, 115]
         16'd223: out = 32'b11010010100000000001111110000000; // MOVZ X0, 252 // Character D
         16'd224: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd225: out = 32'b11110010100111111000000000000000; // MOVK X0, 64512
         16'd226: out = 32'b11111000000001111000001111100000; // STUR X0, [XZR, 120]
         16'd227: out = 32'b11111000000001111100001111100000; // STUR X0, [XZR, 124]
         16'd228: out = 32'b11110010100000000001111110000000; // MOVK X0, 252
         16'd229: out = 32'b11111000000001111001001111100000; // STUR X0, [XZR, 121]
         16'd230: out = 32'b11111000000001111010001111100000; // STUR X0, [XZR, 122]
         16'd231: out = 32'b11111000000001111011001111100000; // STUR X0, [XZR, 123]
         16'd232: out = 32'b11010010100000000001111110000000; // MOVZ X0, 252 // Character E
         16'd233: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd234: out = 32'b11111000000010000001001111100000; // STUR X0, [XZR, 129]
         16'd235: out = 32'b11111000000010000011001111100000; // STUR X0, [XZR, 131]
         16'd236: out = 32'b11110010100111111001111110000000; // MOVK X0, 64764
         16'd237: out = 32'b11111000000010000000001111100000; // STUR X0, [XZR, 128]
         16'd238: out = 32'b11111000000010000100001111100000; // STUR X0, [XZR, 132]
         16'd239: out = 32'b11110010100111111000000000000000; // MOVK X0, 64512
         16'd240: out = 32'b11111000000010000010001111100000; // STUR X0, [XZR, 130]
         16'd241: out = 32'b11010010100000000001111110000000; // MOVZ X0, 252 // Character F
         16'd242: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd243: out = 32'b11111000000010001001001111100000; // STUR X0, [XZR, 137]
         16'd244: out = 32'b11111000000010001011001111100000; // STUR X0, [XZR, 139]
         16'd245: out = 32'b11111000000010001100001111100000; // STUR X0, [XZR, 140]
         16'd246: out = 32'b11110010100111111001111110000000; // MOVK X0, 64764
         16'd247: out = 32'b11111000000010001000001111100000; // STUR X0, [XZR, 136]
         16'd248: out = 32'b11110010100111111000000000000000; // MOVK X0, 64512
         16'd249: out = 32'b11111000000010001010001111100000; // STUR X0, [XZR, 138]
         16'd250: out = 32'b11010010100101011001010110000000; // MOVZ X0, 44204 // Start of alien - 176-185
         16'd251: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd252: out = 32'b11110010100101011001100000000000; // MOVK X0, 44224
         16'd253: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd254: out = 32'b11110010100110000001100000000000; // MOVK X0, 49344
         16'd255: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd256: out = 32'b11110010100101011001010110000000; // MOVK X0, 44204
         16'd257: out = 32'b11111000000010110000001111100000; // STUR X0, [XZR, 176]
         16'd258: out = 32'b11010010100101011001100000000000; // MOVZ X0, 44224
         16'd259: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd260: out = 32'b11110010100110000001100000000000; // MOVK X0, 49344
         16'd261: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd262: out = 32'b11110010100110000001100000000000; // MOVK X0, 49344
         16'd263: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd264: out = 32'b11110010100110000001100000000000; // MOVK X0, 49344
         16'd265: out = 32'b11111000000010110001001111100000; // STUR X0, [XZR, 177]
         16'd266: out = 32'b11111000000010110010001111100000; // STUR X0, [XZR, 178]
         16'd267: out = 32'b11111000000010110011001111100000; // STUR X0, [XZR, 179]
         16'd268: out = 32'b11111000000010110100001111100000; // STUR X0, [XZR, 180]
         16'd269: out = 32'b11111000000010110101001111100000; // STUR X0, [XZR, 181]
         16'd270: out = 32'b11111000000010110110001111100000; // STUR X0, [XZR, 182]
         16'd271: out = 32'b11111000000010110111001111100000; // STUR X0, [XZR, 183]
         16'd272: out = 32'b11010010100101011001100000000000; // MOVZ X0, 44224
         16'd273: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd274: out = 32'b11110010100101011001010110000000; // MOVK X0, 44204
         16'd275: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd276: out = 32'b11110010100101011001010110000000; // MOVK X0, 44204
         16'd277: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd278: out = 32'b11110010100101011001100000000000; // MOVK X0, 44224
         16'd279: out = 32'b11111000000010111000001111100000; // STUR X0, [XZR, 184]
         16'd280: out = 32'b11010010100101011001010110000000; // MOVZ X0, 44204
         16'd281: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd282: out = 32'b11110010100110000001100000000000; // MOVK X0, 49344
         16'd283: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd284: out = 32'b11110010100101011001100000000000; // MOVK X0, 44224
         16'd285: out = 32'b11010011011000000100000000000000; // LSL X0, X0, 16
         16'd286: out = 32'b11110010100110000001010110000000; // MOVK X0, 49324
         16'd287: out = 32'b11111000000010111001001111100000; // STUR X0, [XZR, 185]
         16'd288: out = 32'b00010100000000000000000010001010; // B WaitForVSync // Wait for a vsync to occur
         //
         // DisplayGameBoard: // ***** Display the game board, automatically calls DisplayAliens
         16'd289: out = 32'b11010010100000000011110000000010; // MOVZ X2, 480 // Countdown of 480 addresses for the top of the game board
         16'd290: out = 32'b11111000010000000001001111100000; // LDUR X0, [XZR, 1] // Light blue
         16'd291: out = 32'b11111000010000001010001111100001; // LDUR X1, [XZR, 10] // Top address
         // DGB-Top: // Top of the game board
         16'd292: out = 32'b11111000000000000000000000100000; // STUR X0, [X1, 0]
         16'd293: out = 32'b10010001000000000000010000100001; // ADDI X1, X1, 1
         16'd294: out = 32'b11010001000000000000010001000010; // SUBI X2, X2, 1
         16'd295: out = 32'b10110101111111111111111110000010; // CBNZ X2, DGB-Top // Keep displaying this for each 8 pixel block
         16'd296: out = 32'b11010010100000000000011001000010; // MOVZ X2, 50 // Countdown of 50 addresses for the middle of the game board
         16'd297: out = 32'b11111000010000000010001111100000; // LDUR X0, [XZR, 2] // Dark blue
         16'd298: out = 32'b11111000010000001011001111100001; // LDUR X1, [XZR, 11] // Middle address
         // DGB-Middle: // Middle of the game board
         16'd299: out = 32'b11111000000000000000000000100000; // STUR X0, [X1, 0]
         16'd300: out = 32'b10010001000000000000010000100001; // ADDI X1, X1, 1
         16'd301: out = 32'b11010001000000000000010001000010; // SUBI X2, X2, 1
         16'd302: out = 32'b10110101111111111111111110000010; // CBNZ X2, DGB-Middle // Keep displaying this for each 8 pixel block
         16'd303: out = 32'b11010010100000000000100011000010; // MOVZ X2, 70 // Countdown of 70 addresses for the bottom of the game board
         16'd304: out = 32'b11111000010000000011001111100000; // LDUR X0, [XZR, 3] // Brown
         16'd305: out = 32'b11111000010000001100001111100001; // LDUR X1, [XZR, 12] // Top address
         // DGB-Bottom: // Bottom of the game board
         16'd306: out = 32'b11111000000000000000000000100000; // STUR X0, [X1, 0]
         16'd307: out = 32'b10010001000000000000010000100001; // ADDI X1, X1, 1
         16'd308: out = 32'b11010001000000000000010001000010; // SUBI X2, X2, 1
         16'd309: out = 32'b10110101111111111111111110000010; // CBNZ X2, DGB-Bottom // Keep displaying this for each 8 pixel block
         16'd310: out = 32'b00010100000000000000000000000000; // B DisplayAliens
         //
         // DisplayAliens: // ***** Display the aliens on the game board, automatically calls DisplayGameText
         16'd311: out = 32'b11010010100000000000010000000000; // MOVZ X0, 32 // Counter
         // DA-SingleAlien:
         16'd312: out = 32'b11111000010011000000000000000010; // LDUR X2, [X0, 192] // Get the alien data
         16'd313: out = 32'b11010011010000001111110001000011; // LSR X3, X2, 63
         16'd314: out = 32'b10010010000000000011110001000100; // ANDI X4, X2, 15 // Right char
         16'd315: out = 32'b11010011011000000000110010000100; // LSL X4, X4, 3
         16'd316: out = 32'b10010001000000000101110010000100; // ADDI X4, X4, 23
         16'd317: out = 32'b11010011010000000001000001000101; // LSR X5, X2, 4
         16'd318: out = 32'b10010010000000000011110010100101; // ANDI X5, X5, 15 // Left char
         16'd319: out = 32'b11010011011000000000110010100101; // LSL X5, X5, 3
         16'd320: out = 32'b10010001000000000101110010100101; // ADDI X5, X5, 23
         16'd321: out = 32'b11010011010000000010000001000110; // LSR X6, X2, 8
         16'd322: out = 32'b10010010000000111111110011000110; // ANDI X6, X6, 255 // Y
         16'd323: out = 32'b11010010100000000000000000001000; // MOVZ X8, 0
         16'd324: out = 32'b10110100000000000000000001100110; // CBZ X6, DA-SA-SkipYOffset
         // DA-SA-YOffset:
         16'd325: out = 32'b10010001000000000010100100001000; // ADDI X8, X8, 10
         16'd326: out = 32'b11010001000000000000010011000110; // SUBI X6, X6, 1
         16'd327: out = 32'b10110101111111111111111110100110; // CBNZ X6, DA-SA-YOffset
         // DA-SA-SkipYOffset:
         16'd328: out = 32'b11010011011000000100000001000111; // LSL X7, X2, 16
         16'd329: out = 32'b10010010000000111111110011100111; // ANDI X7, X7, 255 // X
         16'd330: out = 32'b10010001000000000000010011100111; // ADDI X7, X7, 1
         16'd331: out = 32'b10001011000001110000000100001000; // ADD X8, X8, X7 // Get the offset for the gpu
         16'd332: out = 32'b11111000010000001010001111101011; // LDUR X11, [XZR, 10]
         16'd333: out = 32'b10001011000010110000000100001000; // ADD X8, X8, X11
         16'd334: out = 32'b10110100000000000000000111000011; // CBZ X3, DA-SkipAlien // Skip the alien if invalid
         16'd335: out = 32'b11010010100000000000000101000001; // MOVZ X1, 10 // Counter
         // DA-SA-Layer:
         16'd336: out = 32'b10010001000000101011110000101001; // ADDI X9, X1, 175
         16'd337: out = 32'b11111000010000000000000100101010; // LDUR X10, [X9, 0]
         16'd338: out = 32'b11111000010000000000000010001100; // LDUR X12, [X4, 0]
         16'd339: out = 32'b11111000010000000000000010101101; // LDUR X13, [X5, 0]
         16'd340: out = 32'b11010011011000001000000110101101; // LSL X13, X13, 32
         16'd341: out = 32'b10101010000011010000000110001100; // ORR X12, X12, X13
         16'd342: out = 32'b10101010000011000000000101001010; // ORR X10, X10, X12
         16'd343: out = 32'b11111000000000000000000100001010; // STUR X10, [X8, 0]
         16'd344: out = 32'b11010001000000000000010010000100; // SUBI X4, X4, 1
         16'd345: out = 32'b11010001000000000000010010100101; // SUBI X5, X5, 1
         16'd346: out = 32'b11010001000000000010100100001000; // SUBI X8, X8, 10
         16'd347: out = 32'b11010001000000000000010000100001; // SUBI X1, X1, 1
         16'd348: out = 32'b10110101111111111111111001100001; // CBNZ X1, DA-SA-Layer
         // DA-SkipAlien: // Only call this when skipping the alien because it is invalid
         16'd349: out = 32'b11010001000000000000010000000000; // SUBI X0, X0, 1
         16'd350: out = 32'b10110101111111111111101100100000; // CBNZ X0, DA-SingleAlien
         16'd351: out = 32'b00010100000000000000000000000000; // B DisplayGameText
         //
         // DisplayGameText: // ***** Display the text overlaid on the game, automatically calls WaitForVSync
         16'd352: out = 32'b11111000010011111100001111100000; // LDUR X0, [XZR, 252] // Load the current input
         16'd353: out = 32'b11111000010000001100001111100001; // LDUR X1, [XZR, 12] // Ground start location
         16'd354: out = 32'b10010001000000000100000000100001; // ADDI X1, X1, 16 // Offset to lsb
         16'd355: out = 32'b11010010100000000000000010001011; // MOVZ X11, 4 // Counter
         // DGT-DoubleCharInput: // Display the input
         16'd356: out = 32'b10010001000000000000000000000010; // ADDI X2, X0, 0
         16'd357: out = 32'b10010001000000000000000000000011; // ADDI X3, X0, 0
         16'd358: out = 32'b10010010000000000000010001000010; // ANDI X2, X2, 1 // Right side
         16'd359: out = 32'b11010011011000000000110001000010; // LSL X2, X2, 3
         16'd360: out = 32'b10010001000000000100000001000010; // ADDI X2, X2, 16
         16'd361: out = 32'b11010011010000000000010001100011; // LSR X3, X3, 1 // Left side
         16'd362: out = 32'b10010010000000000000010001100011; // ANDI X3, X3, 1
         16'd363: out = 32'b11010011011000000000110001100011; // LSL X3, X3, 3
         16'd364: out = 32'b10010001000000000100000001100011; // ADDI X3, X3, 16
         16'd365: out = 32'b11010010100000000000000010101010; // MOVZ X10, 5 // Counter
         // DGT-DCI-CharLayerInput:
         16'd366: out = 32'b11111000010000000000000000100100; // LDUR X4, [X1, 0] // Get the ground
         16'd367: out = 32'b11111000010000000000001111100101; // LDUR X5, [XZR, 0] // Get the white color
         16'd368: out = 32'b11111000010000000000000001001000; // LDUR X8, [X2, 0] // Get the right char layer
         16'd369: out = 32'b11111000010000000000000001101001; // LDUR X9, [X3, 0] // Get the left char layer
         16'd370: out = 32'b11010011011000001000000100101001; // LSL X9, X9, 32
         16'd371: out = 32'b10001011000010010000000100001000; // ADD X8, X8, X9 // Combine the layers into a bitmask
         16'd372: out = 32'b11001011000010000000001111101001; // SUB X9, XZR, X8
         16'd373: out = 32'b11010001000000000000010100101001; // SUBI X9, X9, 1 // Invert bitmask
         16'd374: out = 32'b10001010000010010000000010000100; // AND X4, X4, X9 // Cut out the new pixels from the background
         16'd375: out = 32'b10001010000010000000000010100101; // AND X5, X5, X8 // Only use the color the bitmask selects
         16'd376: out = 32'b10001011000001010000000010000100; // ADD X4, X4, X5 // Combine the final color in this layer
         16'd377: out = 32'b11111000000000000000000000100100; // STUR X4, [X1, 0] // Store the color
         16'd378: out = 32'b10010001000000000010100000100001; // ADDI X1, X1, 10
         16'd379: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd380: out = 32'b10010001000000000000010001100011; // ADDI X3, X3, 1
         16'd381: out = 32'b11010001000000000000010101001010; // SUBI X10, X10, 1 // Counter
         16'd382: out = 32'b10110101111111111111110111101010; // CBNZ X10, DGT-DCI-CharLayerInput // Display another layer
         16'd383: out = 32'b11010001000000001100110000100001; // SUBI X1, X1, 51
         16'd384: out = 32'b11010011010000000000100000000000; // LSR X0, X0, 2
         16'd385: out = 32'b11010001000000000000010101101011; // SUBI X11, X11, 1 // Counter
         16'd386: out = 32'b10110101111111111111110000101011; // CBNZ X11, DGT-DoubleCharInput // Display another set of characters
         16'd387: out = 32'b11111000010011111010001111100000; // LDUR X0, [XZR, 250] // Load the current score
         16'd388: out = 32'b11111000010000001100001111100001; // LDUR X1, [XZR, 12] // Ground start location
         16'd389: out = 32'b10010001000000000100110000100001; // ADDI X1, X1, 19 // Offset to lsb
         16'd390: out = 32'b11010010100000000000000000101011; // MOVZ X11, 1 // Counter
         // DGT-DoubleCharScore: // Display the score
         16'd391: out = 32'b10010001000000000000000000000010; // ADDI X2, X0, 0
         16'd392: out = 32'b10010001000000000000000000000011; // ADDI X3, X0, 0
         16'd393: out = 32'b10010010000000000011110001000010; // ANDI X2, X2, 15 // Right side
         16'd394: out = 32'b11010011011000000000110001000010; // LSL X2, X2, 3
         16'd395: out = 32'b10010001000000000100000001000010; // ADDI X2, X2, 16
         16'd396: out = 32'b11010011010000000001000001100011; // LSR X3, X3, 4 // Left side
         16'd397: out = 32'b10010010000000000011110001100011; // ANDI X3, X3, 15
         16'd398: out = 32'b11010011011000000000110001100011; // LSL X3, X3, 3
         16'd399: out = 32'b10010001000000000100000001100011; // ADDI X3, X3, 16
         16'd400: out = 32'b11010010100000000000000010101010; // MOVZ X10, 5 // Counter
         // DGT-DCI-CharLayerScore:
         16'd401: out = 32'b11111000010000000000000000100100; // LDUR X4, [X1, 0] // Get the ground
         16'd402: out = 32'b11111000010000000100001111100101; // LDUR X5, [XZR, 4] // Get the yellow color
         16'd403: out = 32'b11111000010000000000000001001000; // LDUR X8, [X2, 0] // Get the right char layer
         16'd404: out = 32'b11111000010000000000000001101001; // LDUR X9, [X3, 0] // Get the left char layer
         16'd405: out = 32'b11010011011000001000000100101001; // LSL X9, X9, 32
         16'd406: out = 32'b10001011000010010000000100001000; // ADD X8, X8, X9 // Combine the layers into a bitmask
         16'd407: out = 32'b11001011000010000000001111101001; // SUB X9, XZR, X8
         16'd408: out = 32'b11010001000000000000010100101001; // SUBI X9, X9, 1 // Invert bitmask
         16'd409: out = 32'b10001010000010010000000010000100; // AND X4, X4, X9 // Cut out the new pixels from the background
         16'd410: out = 32'b10001010000010000000000010100101; // AND X5, X5, X8 // Only use the color the bitmask selects
         16'd411: out = 32'b10001011000001010000000010000100; // ADD X4, X4, X5 // Combine the final color in this layer
         16'd412: out = 32'b11111000000000000000000000100100; // STUR X4, [X1, 0] // Store the color
         16'd413: out = 32'b10010001000000000010100000100001; // ADDI X1, X1, 10
         16'd414: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd415: out = 32'b10010001000000000000010001100011; // ADDI X3, X3, 1
         16'd416: out = 32'b11010001000000000000010101001010; // SUBI X10, X10, 1 // Counter
         16'd417: out = 32'b10110101111111111111110111101010; // CBNZ X10, DGT-DCI-CharLayerScore // Display another layer
         16'd418: out = 32'b11010001000000001100110000100001; // SUBI X1, X1, 51
         16'd419: out = 32'b11010011010000000000100000000000; // LSR X0, X0, 2
         16'd420: out = 32'b11010001000000000000010101101011; // SUBI X11, X11, 1 // Counter
         16'd421: out = 32'b10110101111111111111110000101011; // CBNZ X11, DGT-DoubleCharScore // Display another set of characters
         16'd422: out = 32'b00010100000000000000000000000000; // B UpdateDisplay
         //
         // UpdateDisplay: // ***** Load the pixel data and set into pixel mode
         16'd423: out = 32'b11010010100000000000000010100000; // MOVZ X0, 5 // Set the GPU into pixel and load mode
         16'd424: out = 32'b11111000010000001000001111100001; // LDUR X1, [XZR, 8] // Control address
         16'd425: out = 32'b11111000000000000000000000100000; // STUR X0, [X1, 0]
         16'd426: out = 32'b00010100000000000000000000000000; // B WaitForVSync
         //
         // WaitForVSync: // ***** Wait for the next vsync to pass and CheckForKeyboard, automatically calls DisplayGameBoard
         16'd427: out = 32'b11111000010000001001001111100001; // LDUR X1, [XZR, 9] // Status address for GPU
         // WFVVRise:
         16'd428: out = 32'b10010100000000000000000000010111; // BL CheckForKeyboard // Check for keyboard event and handle it
         16'd429: out = 32'b11111000010000000000000000100000; // LDUR X0, [X1, 0] // Load the status
         16'd430: out = 32'b10010010000000000000100000000000; // ANDI X0, X0, 2
         16'd431: out = 32'b10110100111111111111111110000000; // CBZ X0, WFVVRise // Jump back while vsync is low
         // WFV-DisplayEnableRise:
         16'd432: out = 32'b10010100000000000000000000010011; // BL CheckForKeyboard // Check for keyboard event and handle it
         16'd433: out = 32'b11111000010000000000000000100000; // LDUR X0, [X1, 0] // Load the status
         16'd434: out = 32'b10010010000000000000010000000000; // ANDI X0, X0, 1
         16'd435: out = 32'b10110100111111111111111110000000; // CBZ X0, WFV-DisplayEnableRise // Jump back while display enable is low
         16'd436: out = 32'b00010100000000000000000000000000; // B DoGame
         //
         // DoGame: // ***** Game calcuations
         16'd437: out = 32'b11111000010011111100001111100101; // LDUR X5, [XZR, 252]
         16'd438: out = 32'b11010010100000000000010000000000; // MOVZ X0, 32 // Counter
         // DG-AlienDestroy:
         16'd439: out = 32'b11111000010010111111000000000001; // LDUR X1, [X0, 191]
         16'd440: out = 32'b11010011010000001111110000100010; // LSR X2, X1, 63
         16'd441: out = 32'b10110100000000000000000011100010; // CBZ X2, DG-AD-Skip // Alien already destroyed
         16'd442: out = 32'b10010010000000111111110000100011; // ANDI X3, X1, 255
         16'd443: out = 32'b11001011000001010000000001100100; // SUB X4, X3, X5
         16'd444: out = 32'b10110101000000000000000010000100; // CBNZ X4, DG-AD-Skip // Don't match codes
         16'd445: out = 32'b11111000000010111111000000011111; // STUR XZR, [X0, 191]
         16'd446: out = 32'b11111000010011111010001111100110; // LDUR X6, [XZR, 250]
         16'd447: out = 32'b10010001000000000000010011000110; // ADDI X6, X6, 1
         16'd448: out = 32'b11111000000011111010001111100110; // STUR X6, [XZR, 250]
         // DG-AD-Skip:
         16'd449: out = 32'b11010001000000000000010000000000; // SUBI X0, X0, 1
         16'd450: out = 32'b10110101111111111111111010000000; // CBNZ X0, DG-AlienDestroy
         16'd451: out = 32'b00010111111111111111111101011101; // B DisplayGameBoard
         //
         // CheckForKeyboard: // ***** Check for new keyboard data, if new it calls OnKeyboardPress
         16'd452: out = 32'b10010001000000000000001111011101; // ADDI X29, X30, 0 // Store the location the call came from
         16'd453: out = 32'b11111000010011111110001111110100; // LDUR X20, [XZR, 254] // Get keyboard address
         16'd454: out = 32'b11111000010000000000001010010100; // LDUR X20, [X20, 0] // Get the first keyboard register data
         16'd455: out = 32'b11010011010000000011101010010100; // LSR X20, X20, 14
         16'd456: out = 32'b10010010000000111111111010010100; // ANDI X20, X20, 255 // Isolate the 1-8 keys
         16'd457: out = 32'b10110100000000000000000000110100; // CBZ X20, CFK-NoKeyboard
         16'd458: out = 32'b10010100000000000000000000000010; // BL OnKeyboardPress // Handle keyboard press
         // CFK-NoKeyboard:
         16'd459: out = 32'b11111000000011111101001111110100; // STUR X20, [XZR, 253] // Store the new last keyboard input
         16'd460: out = 32'b11010110000000000000001110100000; // BR X29 // Return to the calling location
         //
         // OnKeyboardPress: // ***** Depending on the state of the game, update the game state
         16'd461: out = 32'b11111000010011111100001111110111; // LDUR X23, [XZR, 252] // Input
         16'd462: out = 32'b11111000010011111101001111111000; // LDUR X24, [XZR, 253] // Last keyboard input
         16'd463: out = 32'b11111000010000000000001111111010; // LDUR X26, [XZR, 0] // White
         16'd464: out = 32'b11111000010000001010001111111011; // LDUR X27, [XZR, 10] // Top of GPU
         16'd465: out = 32'b11001011000110000000001111110101; // SUB X21, XZR, X24
         16'd466: out = 32'b11010001000000000000011010110101; // SUBI X21, X21, 1 // Invert last keyboard
         16'd467: out = 32'b11010011010000000001111010011100; // LSR X28, X20, 7 // Flip the keyboard data bits
         16'd468: out = 32'b10010010000000000000011110011100; // ANDI X28, X28, 1
         16'd469: out = 32'b11010011010000000001011010010011; // LSR X19, X20, 5
         16'd470: out = 32'b10010010000000000000101001110011; // ANDI X19, X19, 2
         16'd471: out = 32'b10101010000100110000001110011100; // ORR X28, X28, X19
         16'd472: out = 32'b11010011010000000000111010010011; // LSR X19, X20, 3
         16'd473: out = 32'b10010010000000000001001001110011; // ANDI X19, X19, 4
         16'd474: out = 32'b10101010000100110000001110011100; // ORR X28, X28, X19
         16'd475: out = 32'b11010011010000000000011010010011; // LSR X19, X20, 1
         16'd476: out = 32'b10010010000000000010001001110011; // ANDI X19, X19, 8
         16'd477: out = 32'b10101010000100110000001110011100; // ORR X28, X28, X19
         16'd478: out = 32'b11010011011000000000011010010011; // LSL X19, X20, 1
         16'd479: out = 32'b10010010000000000100001001110011; // ANDI X19, X19, 16
         16'd480: out = 32'b10101010000100110000001110011100; // ORR X28, X28, X19
         16'd481: out = 32'b11010011011000000000111010010011; // LSL X19, X20, 3
         16'd482: out = 32'b10010010000000001000001001110011; // ANDI X19, X19, 32
         16'd483: out = 32'b10101010000100110000001110011100; // ORR X28, X28, X19
         16'd484: out = 32'b11010011011000000001011010010011; // LSL X19, X20, 5
         16'd485: out = 32'b10010010000000010000001001110011; // ANDI X19, X19, 64
         16'd486: out = 32'b10101010000100110000001110011100; // ORR X28, X28, X19
         16'd487: out = 32'b11010011011000000001111010010011; // LSL X19, X20, 7
         16'd488: out = 32'b10010010000000100000001001110011; // ANDI X19, X19, 128
         16'd489: out = 32'b10101010000100110000001110011100; // ORR X28, X28, X19
         16'd490: out = 32'b10001011000111110000001110010100; // ADD X20, X28, XZR // Copy the keyboard data bits back in
         16'd491: out = 32'b10010010000000000000011010010110; // ANDI X22, X20, 1
         16'd492: out = 32'b10110100000000000000000011010110; // CBZ X22, OKB-Skip1
         16'd493: out = 32'b10010010000000000000011010111001; // ANDI X25, X21, 1
         16'd494: out = 32'b10001010000101100000001100111001; // AND X25, X25, X22
         16'd495: out = 32'b10110100000000000000000001111001; // CBZ X25, OKB-Skip1
         16'd496: out = 32'b11001010000110010000001011110111; // EOR X23, X23, X25
         16'd497: out = 32'b11111000000011111100001111110111; // STUR X23, [XZR, 252]
         16'd498: out = 32'b11010110000000000000001111000000; // BR X30
         // OKB-Skip1:
         16'd499: out = 32'b10010010000000000000101010010110; // ANDI X22, X20, 2
         16'd500: out = 32'b10110100000000000000000011010110; // CBZ X22, OKB-Skip2
         16'd501: out = 32'b10010010000000000000101010111001; // ANDI X25, X21, 2
         16'd502: out = 32'b10001010000101100000001100111001; // AND X25, X25, X22
         16'd503: out = 32'b10110100000000000000000001111001; // CBZ X25, OKB-Skip2
         16'd504: out = 32'b11001010000110010000001011110111; // EOR X23, X23, X25
         16'd505: out = 32'b11111000000011111100001111110111; // STUR X23, [XZR, 252]
         16'd506: out = 32'b11010110000000000000001111000000; // BR X30
         // OKB-Skip2:
         16'd507: out = 32'b10010010000000000001001010010110; // ANDI X22, X20, 4
         16'd508: out = 32'b10110100000000000000000011010110; // CBZ X22, OKB-Skip3
         16'd509: out = 32'b10010010000000000001001010111001; // ANDI X25, X21, 4
         16'd510: out = 32'b10001010000101100000001100111001; // AND X25, X25, X22
         16'd511: out = 32'b10110100000000000000000001111001; // CBZ X25, OKB-Skip3
         16'd512: out = 32'b11001010000110010000001011110111; // EOR X23, X23, X25
         16'd513: out = 32'b11111000000011111100001111110111; // STUR X23, [XZR, 252]
         16'd514: out = 32'b11010110000000000000001111000000; // BR X30
         // OKB-Skip3:
         16'd515: out = 32'b10010010000000000010001010010110; // ANDI X22, X20, 8
         16'd516: out = 32'b10110100000000000000000011010110; // CBZ X22, OKB-Skip4
         16'd517: out = 32'b10010010000000000010001010111001; // ANDI X25, X21, 8
         16'd518: out = 32'b10001010000101100000001100111001; // AND X25, X25, X22
         16'd519: out = 32'b10110100000000000000000001111001; // CBZ X25, OKB-Skip4
         16'd520: out = 32'b11001010000110010000001011110111; // EOR X23, X23, X25
         16'd521: out = 32'b11111000000011111100001111110111; // STUR X23, [XZR, 252]
         16'd522: out = 32'b11010110000000000000001111000000; // BR X30
         // OKB-Skip4:
         16'd523: out = 32'b10010010000000000100001010010110; // ANDI X22, X20, 16
         16'd524: out = 32'b10110100000000000000000011010110; // CBZ X22, OKB-Skip5
         16'd525: out = 32'b10010010000000000100001010111001; // ANDI X25, X21, 16
         16'd526: out = 32'b10001010000101100000001100111001; // AND X25, X25, X22
         16'd527: out = 32'b10110100000000000000000001111001; // CBZ X25, OKB-Skip5
         16'd528: out = 32'b11001010000110010000001011110111; // EOR X23, X23, X25
         16'd529: out = 32'b11111000000011111100001111110111; // STUR X23, [XZR, 252]
         16'd530: out = 32'b11010110000000000000001111000000; // BR X30
         // OKB-Skip5:
         16'd531: out = 32'b10010010000000001000001010010110; // ANDI X22, X20, 32
         16'd532: out = 32'b10110100000000000000000011010110; // CBZ X22, OKB-Skip6
         16'd533: out = 32'b10010010000000001000001010111001; // ANDI X25, X21, 32
         16'd534: out = 32'b10001010000101100000001100111001; // AND X25, X25, X22
         16'd535: out = 32'b10110100000000000000000001111001; // CBZ X25, OKB-Skip6
         16'd536: out = 32'b11001010000110010000001011110111; // EOR X23, X23, X25
         16'd537: out = 32'b11111000000011111100001111110111; // STUR X23, [XZR, 252]
         16'd538: out = 32'b11010110000000000000001111000000; // BR X30
         // OKB-Skip6:
         16'd539: out = 32'b10010010000000010000001010010110; // ANDI X22, X20, 64
         16'd540: out = 32'b10110100000000000000000011010110; // CBZ X22, OKB-Skip7
         16'd541: out = 32'b10010010000000010000001010111001; // ANDI X25, X21, 64
         16'd542: out = 32'b10001010000101100000001100111001; // AND X25, X25, X22
         16'd543: out = 32'b10110100000000000000000001111001; // CBZ X25, OKB-Skip7
         16'd544: out = 32'b11001010000110010000001011110111; // EOR X23, X23, X25
         16'd545: out = 32'b11111000000011111100001111110111; // STUR X23, [XZR, 252]
         16'd546: out = 32'b11010110000000000000001111000000; // BR X30
         // OKB-Skip7:
         16'd547: out = 32'b10010010000000100000001010010110; // ANDI X22, X20, 128
         16'd548: out = 32'b10110100000000000000000011010110; // CBZ X22, OKB-Skip8
         16'd549: out = 32'b10010010000000100000001010111001; // ANDI X25, X21, 128
         16'd550: out = 32'b10001010000101100000001100111001; // AND X25, X25, X22
         16'd551: out = 32'b10110100000000000000000001111001; // CBZ X25, OKB-Skip8
         16'd552: out = 32'b11001010000110010000001011110111; // EOR X23, X23, X25
         16'd553: out = 32'b11111000000011111100001111110111; // STUR X23, [XZR, 252]
         16'd554: out = 32'b11010110000000000000001111000000; // BR X30
         // OKB-Skip8:
         16'd555: out = 32'b11010110000000000000001111000000; // BR X30
         default: out = 32'b11010110000000000000001111100000; // BR XZR
      endcase
   end
endmodule
