module SD_Card;

endmodule
