module ROM_GPIO_Image(out, address);
output reg [31:0] out;
input  [15:0] address; // address- 16 deep memory  
always @(address) begin
case (address)
16'h0000:  out = 32'b11010010100000000000000010100001; // MOVZ X1, 5			// set registry to allocated memory
16'h0001:  out = 32'b11010011011000001110000000100001; // LSL X1, X1, 56
16'h0002:  out = 32'b11010010100000000000000101111101; // MOVZ X29, 11		//store line number
16'h0003:  out = 32'b11110010100100000000000000101010; // MOVK X10, 32769		// load top half of image into register
16'h0004:  out = 32'b11010011011000000100000101001010; // LSL X10, X10, 16
16'h0005:  out = 32'b11110010100100000000000000101010; // MOVK X10, 32769
16'h0006:  out = 32'b11010011011000000100000101001010; // LSL X10, X10, 16
16'h0007:  out = 32'b11110010100100000000000000101010; // MOVK X10, 32769
16'h0008:  out = 32'b11010011011000000100000101001010; // LSL X10, X10, 16
16'h0009:  out = 32'b11110010100100000000000000101010; // MOVK X10, 32769
16'h000a:  out = 32'b11110010100000000000000000010100; // MOVK X20, 0			// load bottom half of image into register
16'h000b:  out = 32'b11010011011000000100001010010100; // LSL X20, X20, 16
16'h000c:  out = 32'b11110010100000000000000000010100; // MOVK X20, 0
16'h000d:  out = 32'b11010011011000000100001010010100; // LSL X20, X20, 16
16'h000e:  out = 32'b11110010100000000000000000010100; // MOVK X20, 0
16'h000f:  out = 32'b11010011011000000100001010010100; // LSL X20, X20, 16
16'h0010:  out = 32'b11110010100000000000000000010100; // MOVK X20, 0
16'h0011:  out = 32'b11111000000000000001000000111111; // STUR XZR, [X1, 1]	// store and load image
16'h0012:  out = 32'b11111000000000000010000000111111; // STUR XZR, [X1, 2]
16'h0013:  out = 32'b11111000000000000011000000111111; // STUR XZR, [X1, 3]
16'h0014:  out = 32'b11111000000000000001000000101010; // STUR X10, [X1, 1]	// store and load image
16'h0015:  out = 32'b11111000000000000010000000110100; // STUR X20, [X1, 2]
16'h0016:  out = 32'b11111000010000000011000000111110; // LDUR X30, [X1, 3]
16'h0017:  out = 32'b11111000000000000011000000111110; // STUR X30, [X1, 3]
16'h0018:  out = 32'b11010010100000000000000000001011; // MOVZ X11, 0
16'h0019:  out = 32'b11010010100000000000000000001101; // MOVZ X13, 0
16'h001a:  out = 32'b11010011011000001100001010001101; // LSL X13, X20, 48	//down
16'h001b:  out = 32'b11010011011000001100000101001011; // LSL X11, X10, 48
16'h001c:  out = 32'b11010011010000000100000101001010; // LSR X10, X10, 16
16'h001d:  out = 32'b11010011010000000100001010010100; // LSR X20, X20, 16
16'h001e:  out = 32'b10001011000011010000000101001010; // ADD X10, X10, X13
16'h001f:  out = 32'b10001011000010110000001010010100; // ADD X20, X20, X11	//end of down
16'h0020:  out = 32'b11111000000000000011000000111111; // STUR XZR, [X1, 3]
16'h0021:  out = 32'b11111000010000000011000000111110; // LDUR X30, [X1, 3]
16'h0022:  out = 32'b11111000000000000011000000111110; // STUR X30, [X1, 3]
16'h0023:  out = 32'b11110001000000000100001111000010; // SUBIS X2, X30, 16
16'h0024:  out = 32'b01010100111111111111111110000001; // B.NE -4			//branch to line 17
16'h0025:  out = 32'b11111000000000000011000000111111; // STUR XZR, [X1, 3]
16'h0026:  out = 32'b11111000010000000011000000111110; // LDUR X30, [X1, 3]
16'h0027:  out = 32'b11111000000000000011000000111110; // STUR X30, [X1, 3]
16'h0028:  out = 32'b11110001000000000100001111000010; // SUBIS X2, X30, 16
16'h0029:  out = 32'b01010100111111111111111110000000; // B.EQ -4
16'h002a:  out = 32'b01010100111111111111110011100001; // B.NE -25
default: out=32'hD60003E0; //BR XZR
endcase
end
endmodule
