module SD_Card(clock, command, data, write_protect);
input clock, write_protect;
inout command, data[1:0];



endmodule
