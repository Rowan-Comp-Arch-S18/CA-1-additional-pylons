module SD_Card(clock, command, data, write_protect);
input write_protect;
output clock;
inout command;
inout [1:0]data;



endmodule
