module ROM_Image_Display(out, address);
   input[15:0] address;
   output reg[31:0] out;
   always @(address) begin
      case(address)
         16'd0: out = 32'b11010010100000000000000001010100; // MOVZ X20, 2
         16'd1: out = 32'b11010011011000001110001010010100; // LSL X20, X20, 56
         16'd2: out = 32'b10010001000000000000101010010101; // ADDI X21, X20, 2
         16'd3: out = 32'b10010001000010010111001010010110; // ADDI X22, X20, 604
         16'd4: out = 32'b10001011000111110000001011000010; // ADD X2, X22, XZR
         16'd5: out = 32'b11111000010000000000001010100011; // LDUR X3, [X21, 0]
         16'd6: out = 32'b10010010000000000000100001100011; // ANDI X3, X3, 2
         16'd7: out = 32'b10110100111111111111111110100011; // CBZ X3, -3
         16'd8: out = 32'b11111000010000000000001010100011; // LDUR X3, [X21, 0]
         16'd9: out = 32'b10010010000000000000010001100011; // ANDI X3, X3, 1
         16'd10: out = 32'b10110100111111111111111110100011; // CBZ X3, -3
         16'd11: out = 32'b11010010100010100000101000000101; // MOVZ X5, 20560
         16'd12: out = 32'b10001011000010100000000010101010; // ADD X10, X5, X10
         16'd13: out = 32'b11010011011000000100000010100101; // LSL X5, X5, 16
         16'd14: out = 32'b10001011000010100000000010101010; // ADD X10, X5, X10
         16'd15: out = 32'b11010011011000000100000010100101; // LSL X5, X5, 16
         16'd16: out = 32'b10001011000010100000000010101010; // ADD X10, X5, X10
         16'd17: out = 32'b11010011011000000100000010100101; // LSL X5, X5, 16
         16'd18: out = 32'b10001011000010100000000010101010; // ADD X10, X5, X10
         16'd19: out = 32'b11010010100111001010001100000110; // MOVZ X6, 58648
         16'd20: out = 32'b10001011000010110000000011001011; // ADD X11, X6, X11
         16'd21: out = 32'b11010011011000000100000011000110; // LSL X6, X6, 16
         16'd22: out = 32'b10001011000010110000000011001011; // ADD X11, X6, X11
         16'd23: out = 32'b11010011011000000100000011000110; // LSL X6, X6, 16
         16'd24: out = 32'b10001011000010110000000011001011; // ADD X11, X6, X11
         16'd25: out = 32'b11010011011000000100000011000110; // LSL X6, X6, 16
         16'd26: out = 32'b10001011000010110000000011001011; // ADD X11, X6, X11
         16'd27: out = 32'b11010010100010101000101010000111; // MOVZ X7, 21588
         16'd28: out = 32'b10001011000011000000000011101100; // ADD X12, X7, X12
         16'd29: out = 32'b11010011011000000100000011100111; // LSL X7, X7, 16
         16'd30: out = 32'b10001011000011000000000011101100; // ADD X12, X7, X12
         16'd31: out = 32'b11010011011000000100000011100111; // LSL X7, X7, 16
         16'd32: out = 32'b10001011000011000000000011101100; // ADD X12, X7, X12
         16'd33: out = 32'b11010011011000000100000011100111; // LSL X7, X7, 16
         16'd34: out = 32'b10001011000011000000000011101100; // ADD X12, X7, X12
         16'd35: out = 32'b11010010100111110001111100001000; // MOVZ X8, 63736
         16'd36: out = 32'b10001011000011010000000100001101; // ADD X13, X8, X13
         16'd37: out = 32'b11010011011000000100000100001000; // LSL X8, X8, 16
         16'd38: out = 32'b10001011000011010000000100001101; // ADD X13, X8, X13
         16'd39: out = 32'b11010011011000000100000100001000; // LSL X8, X8, 16
         16'd40: out = 32'b10001011000011010000000100001101; // ADD X13, X8, X13
         16'd41: out = 32'b11010011011000000100000100001000; // LSL X8, X8, 16
         16'd42: out = 32'b10001011000011010000000100001101; // ADD X13, X8, X13
         16'd43: out = 32'b11010010100111111001111110001001; // MOVZ X9, 64764
         16'd44: out = 32'b10001011000011100000000100101110; // ADD X14, X9, X14
         16'd45: out = 32'b11010011011000000100000100101001; // LSL X9, X9, 16
         16'd46: out = 32'b10001011000011100000000100101110; // ADD X14, X9, X14
         16'd47: out = 32'b11010011011000000100000100101001; // LSL X9, X9, 16
         16'd48: out = 32'b10001011000011100000000100101110; // ADD X14, X9, X14
         16'd49: out = 32'b11010011011000000100000100101001; // LSL X9, X9, 16
         16'd50: out = 32'b10001011000011100000000100101110; // ADD X14, X9, X14
         16'd51: out = 32'b11010010100011001000110010001001; // MOVZ X9, 25700
         16'd52: out = 32'b10001011000011110000000100101111; // ADD X15, X9, X15
         16'd53: out = 32'b11010011011000000100000100101001; // LSL X9, X9, 16
         16'd54: out = 32'b10001011000011110000000100101111; // ADD X15, X9, X15
         16'd55: out = 32'b11010011011000000100000100101001; // LSL X9, X9, 16
         16'd56: out = 32'b10001011000011110000000100101111; // ADD X15, X9, X15
         16'd57: out = 32'b11010011011000000100000100101001; // LSL X9, X9, 16
         16'd58: out = 32'b10001011000011110000000100101111; // ADD X15, X9, X15
         16'd59: out = 32'b11010010100101001001010010001001; // MOVZ X9, 42148
         16'd60: out = 32'b10001011000100000000000100110000; // ADD X16, X9, X16
         16'd61: out = 32'b11010011011000000100000100101001; // LSL X9, X9, 16
         16'd62: out = 32'b10001011000100000000000100110000; // ADD X16, X9, X16
         16'd63: out = 32'b11010011011000000100000100101001; // LSL X9, X9, 16
         16'd64: out = 32'b10001011000100000000000100110000; // ADD X16, X9, X16
         16'd65: out = 32'b11010011011000000100000100101001; // LSL X9, X9, 16
         16'd66: out = 32'b10001011000100000000000100110000; // ADD X16, X9, X16
         16'd67: out = 32'b11010010100111010001110100001001; // MOVZ X9, 59624
         16'd68: out = 32'b10001011000100010000000100110001; // ADD X17, X9, X17
         16'd69: out = 32'b11010011011000000100000100101001; // LSL X9, X9, 16
         16'd70: out = 32'b10001011000100010000000100110001; // ADD X17, X9, X17
         16'd71: out = 32'b11010011011000000100000100101001; // LSL X9, X9, 16
         16'd72: out = 32'b10001011000100010000000100110001; // ADD X17, X9, X17
         16'd73: out = 32'b11010011011000000100000100101001; // LSL X9, X9, 16
         16'd74: out = 32'b10001011000100010000000100110001; // ADD X17, X9, X17
         16'd75: out = 32'b11010010100000001000000010001001; // MOVZ X9, 1028
         16'd76: out = 32'b10001011000100110000000100110011; // ADD X19, X9, X19
         16'd77: out = 32'b11010011011000000100000100101001; // LSL X9, X9, 16
         16'd78: out = 32'b10001011000100110000000100110011; // ADD X19, X9, X19
         16'd79: out = 32'b11010011011000000100000100101001; // LSL X9, X9, 16
         16'd80: out = 32'b10001011000100110000000100110011; // ADD X19, X9, X19
         16'd81: out = 32'b11010011011000000100000100101001; // LSL X9, X9, 16
         16'd82: out = 32'b10001011000100110000000100110011; // ADD X19, X9, X19
         16'd83: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd84: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd85: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd86: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd87: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd88: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd89: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd90: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd91: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd92: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd93: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd94: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd95: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd96: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd97: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd98: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd99: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd100: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd101: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd102: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd103: out = 32'b11110010100000000000000010000001; // MOVK X1, 4
         16'd104: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd105: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd106: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd107: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd108: out = 32'b11010010100010001000101010000001; // MOVZ X1, 17492
         16'd109: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd110: out = 32'b11110010100010101000101010000001; // MOVK X1, 21588
         16'd111: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd112: out = 32'b11110010100010101000101010000001; // MOVK X1, 21588
         16'd113: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd114: out = 32'b11110010100010101000101010000001; // MOVK X1, 21588
         16'd115: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd116: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd117: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd118: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd119: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd120: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd121: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd122: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd123: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd124: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd125: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd126: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd127: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd128: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd129: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd130: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd131: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd132: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd133: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd134: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd135: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd136: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd137: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd138: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd139: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd140: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd141: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd142: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd143: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd144: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd145: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd146: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd147: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd148: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd149: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd150: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd151: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd152: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd153: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd154: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd155: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd156: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd157: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd158: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd159: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd160: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd161: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd162: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd163: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd164: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd165: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd166: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd167: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd168: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd169: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd170: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd171: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd172: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd173: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd174: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd175: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd176: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd177: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd178: out = 32'b11110010100000000000100010000001; // MOVK X1, 68
         16'd179: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd180: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd181: out = 32'b11010010100010101000100000000001; // MOVZ X1, 21568
         16'd182: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd183: out = 32'b11110010100010000000101010000001; // MOVK X1, 16468
         16'd184: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd185: out = 32'b11110010100010101000101010000001; // MOVK X1, 21588
         16'd186: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd187: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd188: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd189: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd190: out = 32'b11010010100010000000000000000001; // MOVZ X1, 16384
         16'd191: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd192: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd193: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd194: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd195: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd196: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd197: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd198: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd199: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd200: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd201: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd202: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd203: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd204: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd205: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd206: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd207: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd208: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd209: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd210: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd211: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd212: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd213: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd214: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd215: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd216: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd217: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd218: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd219: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd220: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd221: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd222: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd223: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd224: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd225: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd226: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd227: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd228: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd229: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd230: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd231: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd232: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd233: out = 32'b11110010100010001000101010000001; // MOVK X1, 17492
         16'd234: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd235: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd236: out = 32'b11010010100010100000101000000001; // MOVZ X1, 20560
         16'd237: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd238: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd239: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd240: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd241: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd242: out = 32'b11110010100010100000101010000001; // MOVK X1, 20564
         16'd243: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd244: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd245: out = 32'b11010010100010100000100000000001; // MOVZ X1, 20544
         16'd246: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd247: out = 32'b11110010100010101000101000000001; // MOVK X1, 21584
         16'd248: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd249: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd250: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd251: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd252: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd253: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd254: out = 32'b11010010100000000000000010000001; // MOVZ X1, 4
         16'd255: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd256: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd257: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd258: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd259: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd260: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd261: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd262: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd263: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd264: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd265: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd266: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd267: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd268: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd269: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd270: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd271: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd272: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd273: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd274: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd275: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd276: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd277: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd278: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd279: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd280: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd281: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd282: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd283: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd284: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd285: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd286: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd287: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd288: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd289: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd290: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd291: out = 32'b11010010100010000000100000000001; // MOVZ X1, 16448
         16'd292: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd293: out = 32'b11110010100010100000101010000001; // MOVK X1, 20564
         16'd294: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd295: out = 32'b11110010100010101000101010000001; // MOVK X1, 21588
         16'd296: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd297: out = 32'b11110010100010101000100000000001; // MOVK X1, 21568
         16'd298: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd299: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd300: out = 32'b11010010100000000000100000000001; // MOVZ X1, 64
         16'd301: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd302: out = 32'b11110010100010101001010010000001; // MOVK X1, 21668
         16'd303: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd304: out = 32'b11110010100010101000000000000001; // MOVK X1, 21504
         16'd305: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd306: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd307: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd308: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd309: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd310: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd311: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd312: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd313: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd314: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd315: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd316: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd317: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd318: out = 32'b11111000000000000000000001010011; // STUR X19, [X2, 0]
         16'd319: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd320: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd321: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd322: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd323: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd324: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd325: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd326: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd327: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd328: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd329: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd330: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd331: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd332: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd333: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd334: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd335: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd336: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd337: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd338: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd339: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd340: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd341: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd342: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd343: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd344: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd345: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd346: out = 32'b11010010100000000000100000000001; // MOVZ X1, 64
         16'd347: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd348: out = 32'b11110010100010101001001010000001; // MOVK X1, 21652
         16'd349: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd350: out = 32'b11110010100100101001010100000001; // MOVK X1, 38056
         16'd351: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd352: out = 32'b11110010100101001000101010000001; // MOVK X1, 42068
         16'd353: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd354: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd355: out = 32'b11010010100010000000100000000001; // MOVZ X1, 16448
         16'd356: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd357: out = 32'b11110010100010000000101010000001; // MOVK X1, 16468
         16'd358: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd359: out = 32'b11110010100010101000000000000001; // MOVK X1, 21504
         16'd360: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd361: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd362: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd363: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd364: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd365: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd366: out = 32'b11110010100000000000000010000001; // MOVK X1, 4
         16'd367: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd368: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd369: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd370: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd371: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd372: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd373: out = 32'b11111000000000000000000001010011; // STUR X19, [X2, 0]
         16'd374: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd375: out = 32'b11111000000000000000000001010011; // STUR X19, [X2, 0]
         16'd376: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd377: out = 32'b11111000000000000000000001010011; // STUR X19, [X2, 0]
         16'd378: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd379: out = 32'b11010010100000001000000000000001; // MOVZ X1, 1024
         16'd380: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd381: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd382: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd383: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd384: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd385: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd386: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd387: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd388: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd389: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd390: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd391: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd392: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd393: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd394: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd395: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd396: out = 32'b11110010100000000000100000000001; // MOVK X1, 64
         16'd397: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd398: out = 32'b11110010100010101001010010000001; // MOVK X1, 21668
         16'd399: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd400: out = 32'b11110010100111010001010100000001; // MOVK X1, 59560
         16'd401: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd402: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd403: out = 32'b11010010100100101000101000000001; // MOVZ X1, 37968
         16'd404: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd405: out = 32'b11110010100010101000101010000001; // MOVK X1, 21588
         16'd406: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd407: out = 32'b11110010100010101000000000000001; // MOVK X1, 21504
         16'd408: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd409: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd410: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd411: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd412: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd413: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd414: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd415: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd416: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd417: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd418: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd419: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd420: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd421: out = 32'b11111000000000000000000001010011; // STUR X19, [X2, 0]
         16'd422: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd423: out = 32'b11111000000000000000000001010011; // STUR X19, [X2, 0]
         16'd424: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd425: out = 32'b11111000000000000000000001010011; // STUR X19, [X2, 0]
         16'd426: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd427: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd428: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd429: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd430: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd431: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd432: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd433: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd434: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd435: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd436: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd437: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd438: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd439: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd440: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd441: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd442: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd443: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd444: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd445: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd446: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd447: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd448: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd449: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd450: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd451: out = 32'b11110010100000000000100000000001; // MOVK X1, 64
         16'd452: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd453: out = 32'b11110010100010100001001010000001; // MOVK X1, 20628
         16'd454: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd455: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd456: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd457: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd458: out = 32'b11010010100111010001001010000001; // MOVZ X1, 59540
         16'd459: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd460: out = 32'b11110010100010101000101010000001; // MOVK X1, 21588
         16'd461: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd462: out = 32'b11110010100010101000100000000001; // MOVK X1, 21568
         16'd463: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd464: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd465: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd466: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd467: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd468: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd469: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd470: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd471: out = 32'b11110010100000000000000010000001; // MOVK X1, 4
         16'd472: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd473: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd474: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd475: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd476: out = 32'b11111000000000000000000001010011; // STUR X19, [X2, 0]
         16'd477: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd478: out = 32'b11111000000000000000000001010011; // STUR X19, [X2, 0]
         16'd479: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd480: out = 32'b11111000000000000000000001010011; // STUR X19, [X2, 0]
         16'd481: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd482: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd483: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd484: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd485: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd486: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd487: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd488: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd489: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd490: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd491: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd492: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd493: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd494: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd495: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd496: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd497: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd498: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd499: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd500: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd501: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd502: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd503: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd504: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd505: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd506: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd507: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd508: out = 32'b11110010100010000000101010000001; // MOVK X1, 16468
         16'd509: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd510: out = 32'b11110010100100101001110100000001; // MOVK X1, 38120
         16'd511: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd512: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd513: out = 32'b11010010100111010001110100000001; // MOVZ X1, 59624
         16'd514: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd515: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd516: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd517: out = 32'b11110010100010101000100000000001; // MOVK X1, 21568
         16'd518: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd519: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd520: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd521: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd522: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd523: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd524: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd525: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd526: out = 32'b11110010100000000000000010000001; // MOVK X1, 4
         16'd527: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd528: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd529: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd530: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd531: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd532: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd533: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd534: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd535: out = 32'b11110010100010001000000010000001; // MOVK X1, 17412
         16'd536: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd537: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd538: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd539: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd540: out = 32'b11111000000000000000000001010011; // STUR X19, [X2, 0]
         16'd541: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd542: out = 32'b11111000000000000000000001010011; // STUR X19, [X2, 0]
         16'd543: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd544: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd545: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd546: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd547: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd548: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd549: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd550: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd551: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd552: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd553: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd554: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd555: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd556: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd557: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd558: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd559: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd560: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd561: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd562: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd563: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd564: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd565: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd566: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd567: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd568: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd569: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd570: out = 32'b11110010100000000000100000000001; // MOVK X1, 64
         16'd571: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd572: out = 32'b11110010100010000001001010000001; // MOVK X1, 16532
         16'd573: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd574: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd575: out = 32'b11010010100111010001111100000001; // MOVZ X1, 59640
         16'd576: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd577: out = 32'b11110010100111010001010010000001; // MOVK X1, 59556
         16'd578: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd579: out = 32'b11110010100010101000100000000001; // MOVK X1, 21568
         16'd580: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd581: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd582: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd583: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd584: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd585: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd586: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd587: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd588: out = 32'b11110010100000000000000010000001; // MOVK X1, 4
         16'd589: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd590: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd591: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd592: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd593: out = 32'b11111000000000000000000001010011; // STUR X19, [X2, 0]
         16'd594: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd595: out = 32'b11111000000000000000000001010011; // STUR X19, [X2, 0]
         16'd596: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd597: out = 32'b11111000000000000000000001010011; // STUR X19, [X2, 0]
         16'd598: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd599: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd600: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd601: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd602: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd603: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd604: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd605: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd606: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd607: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd608: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd609: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd610: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd611: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd612: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd613: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd614: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd615: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd616: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd617: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd618: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd619: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd620: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd621: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd622: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd623: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd624: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd625: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd626: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd627: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd628: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd629: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd630: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd631: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd632: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd633: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd634: out = 32'b11110010100010000000101000000001; // MOVK X1, 16464
         16'd635: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd636: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd637: out = 32'b11010010100100101001110100000001; // MOVZ X1, 38120
         16'd638: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd639: out = 32'b11110010100111010001010010000001; // MOVK X1, 59556
         16'd640: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd641: out = 32'b11110010100010101000100000000001; // MOVK X1, 21568
         16'd642: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd643: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd644: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd645: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd646: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd647: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd648: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd649: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd650: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd651: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd652: out = 32'b11111000000000000000000001010011; // STUR X19, [X2, 0]
         16'd653: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd654: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd655: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd656: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd657: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd658: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd659: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd660: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd661: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd662: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd663: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd664: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd665: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd666: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd667: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd668: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd669: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd670: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd671: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd672: out = 32'b11010010100000001000000100000001; // MOVZ X1, 1032
         16'd673: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd674: out = 32'b11110010100000010000000010000001; // MOVK X1, 2052
         16'd675: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd676: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd677: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd678: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd679: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd680: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd681: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd682: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd683: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd684: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd685: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd686: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd687: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd688: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd689: out = 32'b11110010100010000000101000000001; // MOVK X1, 16464
         16'd690: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd691: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd692: out = 32'b11010010100100101001110100000001; // MOVZ X1, 38120
         16'd693: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd694: out = 32'b11110010100111010001001010000001; // MOVK X1, 59540
         16'd695: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd696: out = 32'b11110010100010101000100000000001; // MOVK X1, 21568
         16'd697: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd698: out = 32'b11110010100010000000000000000001; // MOVK X1, 16384
         16'd699: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd700: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd701: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd702: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd703: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd704: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd705: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd706: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd707: out = 32'b11010010100000010000000100000001; // MOVZ X1, 2056
         16'd708: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd709: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd710: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd711: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd712: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd713: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd714: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd715: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd716: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd717: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd718: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd719: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd720: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd721: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd722: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd723: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd724: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd725: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd726: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd727: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd728: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd729: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd730: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd731: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd732: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd733: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd734: out = 32'b11010010100000010000000100000001; // MOVZ X1, 2056
         16'd735: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd736: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd737: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd738: out = 32'b11110010100010110000000010000001; // MOVK X1, 22532
         16'd739: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd740: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd741: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd742: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd743: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd744: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd745: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd746: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd747: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd748: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd749: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd750: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd751: out = 32'b11110010100000000000100000000001; // MOVK X1, 64
         16'd752: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd753: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd754: out = 32'b11010010100010101001010100000001; // MOVZ X1, 21672
         16'd755: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd756: out = 32'b11110010100111110001110100000001; // MOVK X1, 63720
         16'd757: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd758: out = 32'b11110010100101001000101010000001; // MOVK X1, 42068
         16'd759: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd760: out = 32'b11110010100010000000000000000001; // MOVK X1, 16384
         16'd761: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd762: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd763: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd764: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd765: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd766: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd767: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd768: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd769: out = 32'b11010010100000010000000100000001; // MOVZ X1, 2056
         16'd770: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd771: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd772: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd773: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd774: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd775: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd776: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd777: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd778: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd779: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd780: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd781: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd782: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd783: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd784: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd785: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd786: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd787: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd788: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd789: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd790: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd791: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd792: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd793: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd794: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd795: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd796: out = 32'b11010010100000010000000100000001; // MOVZ X1, 2056
         16'd797: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd798: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd799: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd800: out = 32'b11110010100010110000000010000001; // MOVK X1, 22532
         16'd801: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd802: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd803: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd804: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd805: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd806: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd807: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd808: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd809: out = 32'b11010010100010000001001010000001; // MOVZ X1, 16532
         16'd810: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd811: out = 32'b11110010100101010001110100000001; // MOVK X1, 43240
         16'd812: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd813: out = 32'b11110010100101001001001010000001; // MOVK X1, 42132
         16'd814: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd815: out = 32'b11110010100010100000100000000001; // MOVK X1, 20544
         16'd816: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd817: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd818: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd819: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd820: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd821: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd822: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd823: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd824: out = 32'b11110010100010101001010100000001; // MOVK X1, 21672
         16'd825: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd826: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd827: out = 32'b11010010100101010001010100000001; // MOVZ X1, 43176
         16'd828: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd829: out = 32'b11110010100101010001010100000001; // MOVK X1, 43176
         16'd830: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd831: out = 32'b11110010100101010000101100000001; // MOVK X1, 43096
         16'd832: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd833: out = 32'b11110010100010110000101010000001; // MOVK X1, 22612
         16'd834: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd835: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd836: out = 32'b11010010100010101000101010000001; // MOVZ X1, 21588
         16'd837: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd838: out = 32'b11110010100010101000101010000001; // MOVK X1, 21588
         16'd839: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd840: out = 32'b11110010100010101000001010000001; // MOVK X1, 21524
         16'd841: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd842: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd843: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd844: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd845: out = 32'b11010010100000010000000100000001; // MOVZ X1, 2056
         16'd846: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd847: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd848: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd849: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd850: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd851: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd852: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd853: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd854: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd855: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd856: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd857: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd858: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd859: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd860: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd861: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd862: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd863: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd864: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd865: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd866: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd867: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd868: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd869: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd870: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd871: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd872: out = 32'b11010010100000010000000100000001; // MOVZ X1, 2056
         16'd873: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd874: out = 32'b11110010100000110000101100000001; // MOVK X1, 6232
         16'd875: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd876: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd877: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd878: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd879: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd880: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd881: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd882: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd883: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd884: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd885: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd886: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd887: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd888: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd889: out = 32'b11110010100000000000100000000001; // MOVK X1, 64
         16'd890: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd891: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd892: out = 32'b11010010100010000000101000000001; // MOVZ X1, 16464
         16'd893: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd894: out = 32'b11110010100100101001010100000001; // MOVK X1, 38056
         16'd895: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd896: out = 32'b11110010100101001001001010000001; // MOVK X1, 42132
         16'd897: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd898: out = 32'b11110010100100101000101000000001; // MOVK X1, 37968
         16'd899: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd900: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd901: out = 32'b11010010100010100000100000000001; // MOVZ X1, 20544
         16'd902: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd903: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd904: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd905: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd906: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd907: out = 32'b11110010100010101001111110000001; // MOVK X1, 21756
         16'd908: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd909: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd910: out = 32'b11111000000000000000000001001110; // STUR X14, [X2, 0]
         16'd911: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd912: out = 32'b11111000000000000000000001001110; // STUR X14, [X2, 0]
         16'd913: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd914: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd915: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd916: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd917: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd918: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd919: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd920: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd921: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd922: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd923: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd924: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd925: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd926: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd927: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd928: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd929: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd930: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd931: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd932: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd933: out = 32'b11010010100000010000000100000001; // MOVZ X1, 2056
         16'd934: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd935: out = 32'b11110010100000010000101100000001; // MOVK X1, 2136
         16'd936: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd937: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd938: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd939: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd940: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd941: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd942: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd943: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd944: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd945: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd946: out = 32'b11010010100000000000100000000001; // MOVZ X1, 64
         16'd947: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd948: out = 32'b11110010100100101001010010000001; // MOVK X1, 38052
         16'd949: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd950: out = 32'b11110010100111010001110010000001; // MOVK X1, 59620
         16'd951: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd952: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd953: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd954: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd955: out = 32'b11010010100100101000101010000001; // MOVZ X1, 37972
         16'd956: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd957: out = 32'b11110010100010000000000000000001; // MOVK X1, 16384
         16'd958: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd959: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd960: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd961: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd962: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd963: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd964: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd965: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd966: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd967: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd968: out = 32'b11110010100000000000101010000001; // MOVK X1, 84
         16'd969: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd970: out = 32'b11110010100010101000101010000001; // MOVK X1, 21588
         16'd971: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd972: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd973: out = 32'b11010010100010101000101010000001; // MOVZ X1, 21588
         16'd974: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd975: out = 32'b11110010100010101000101010000001; // MOVK X1, 21588
         16'd976: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd977: out = 32'b11110010100010110001010100000001; // MOVK X1, 22696
         16'd978: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd979: out = 32'b11110010100101010001010100000001; // MOVK X1, 43176
         16'd980: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd981: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd982: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd983: out = 32'b11010010100000010000000010000001; // MOVZ X1, 2052
         16'd984: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd985: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd986: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd987: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd988: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd989: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd990: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd991: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd992: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd993: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd994: out = 32'b11110010100000000000000010000001; // MOVK X1, 4
         16'd995: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd996: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd997: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd998: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd999: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1000: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1001: out = 32'b11010010100000010000000100000001; // MOVZ X1, 2056
         16'd1002: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1003: out = 32'b11110010100000010000000010000001; // MOVK X1, 2052
         16'd1004: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1005: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd1006: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1007: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1008: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1009: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1010: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1011: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1012: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1013: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1014: out = 32'b11010010100010000000100000000001; // MOVZ X1, 16448
         16'd1015: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1016: out = 32'b11110010100010100001001010000001; // MOVK X1, 20628
         16'd1017: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1018: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd1019: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1020: out = 32'b11110010100100101001010010000001; // MOVK X1, 38052
         16'd1021: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1022: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1023: out = 32'b11010010100111001001010010000001; // MOVZ X1, 58532
         16'd1024: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1025: out = 32'b11110010100010101000000000000001; // MOVK X1, 21504
         16'd1026: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1027: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1028: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1029: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1030: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1031: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1032: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1033: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1034: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1035: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1036: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1037: out = 32'b11010010100000010000000100000001; // MOVZ X1, 2056
         16'd1038: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1039: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1040: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1041: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1042: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1043: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1044: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1045: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1046: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd1047: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1048: out = 32'b11110010100000000000000010000001; // MOVK X1, 4
         16'd1049: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1050: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1051: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1052: out = 32'b11110010100000001000000100000001; // MOVK X1, 1032
         16'd1053: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1054: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1055: out = 32'b11010010100010110000101100000001; // MOVZ X1, 22616
         16'd1056: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1057: out = 32'b11110010100010110000101100000001; // MOVK X1, 22616
         16'd1058: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1059: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd1060: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1061: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1062: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1063: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1064: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1065: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1066: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1067: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1068: out = 32'b11010010100010000000100000000001; // MOVZ X1, 16448
         16'd1069: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1070: out = 32'b11110010100100101001010100000001; // MOVK X1, 38056
         16'd1071: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1072: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd1073: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1074: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd1075: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1076: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1077: out = 32'b11010010100111010001110100000001; // MOVZ X1, 59624
         16'd1078: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1079: out = 32'b11110010100100101000100000000001; // MOVK X1, 37952
         16'd1080: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1081: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1082: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1083: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1084: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1085: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1086: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1087: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1088: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1089: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1090: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1091: out = 32'b11010010100000010000000100000001; // MOVZ X1, 2056
         16'd1092: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1093: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1094: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1095: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd1096: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1097: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1098: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1099: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1100: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd1101: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1102: out = 32'b11110010100000000000000010000001; // MOVK X1, 4
         16'd1103: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1104: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1105: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1106: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd1107: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1108: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1109: out = 32'b11010010100010110000101100000001; // MOVZ X1, 22616
         16'd1110: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1111: out = 32'b11110010100010110000101100000001; // MOVK X1, 22616
         16'd1112: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1113: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd1114: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1115: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1116: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1117: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1118: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1119: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1120: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd1121: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1122: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1123: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1124: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd1125: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1126: out = 32'b11110010100010000000101010000001; // MOVK X1, 16468
         16'd1127: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1128: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1129: out = 32'b11010010100100101001110100000001; // MOVZ X1, 38120
         16'd1130: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1131: out = 32'b11110010100111010001111110000001; // MOVK X1, 59644
         16'd1132: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1133: out = 32'b11110010100111111001111110000001; // MOVK X1, 64764
         16'd1134: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1135: out = 32'b11110010100111110001111100000001; // MOVK X1, 63736
         16'd1136: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1137: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1138: out = 32'b11010010100111010001110100000001; // MOVZ X1, 59624
         16'd1139: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1140: out = 32'b11110010100101001000100000000001; // MOVK X1, 42048
         16'd1141: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1142: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1143: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1144: out = 32'b11110010100010000001001010000001; // MOVK X1, 16532
         16'd1145: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1146: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1147: out = 32'b11010010100100101000101010000001; // MOVZ X1, 37972
         16'd1148: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1149: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1150: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1151: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1152: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1153: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1154: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1155: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1156: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1157: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1158: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1159: out = 32'b11010010100000010000000100000001; // MOVZ X1, 2056
         16'd1160: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1161: out = 32'b11110010100000010000000010000001; // MOVK X1, 2052
         16'd1162: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1163: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd1164: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1165: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1166: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1167: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1168: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd1169: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1170: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1171: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1172: out = 32'b11110010100000001000000100000001; // MOVK X1, 1032
         16'd1173: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1174: out = 32'b11110010100000110000101100000001; // MOVK X1, 6232
         16'd1175: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1176: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1177: out = 32'b11010010100010110000101100000001; // MOVZ X1, 22616
         16'd1178: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1179: out = 32'b11110010100010110000001100000001; // MOVK X1, 22552
         16'd1180: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1181: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1182: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1183: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1184: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1185: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1186: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1187: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1188: out = 32'b11010010100000000000100000000001; // MOVZ X1, 64
         16'd1189: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1190: out = 32'b11110010100010101001001010000001; // MOVK X1, 21652
         16'd1191: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1192: out = 32'b11110010100101001001110100000001; // MOVK X1, 42216
         16'd1193: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1194: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd1195: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1196: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1197: out = 32'b11010010100111110001111110000001; // MOVZ X1, 63740
         16'd1198: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1199: out = 32'b11110010100111111001111110000001; // MOVK X1, 64764
         16'd1200: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1201: out = 32'b11110010100111111001111100000001; // MOVK X1, 64760
         16'd1202: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1203: out = 32'b11110010100111110001110100000001; // MOVK X1, 63720
         16'd1204: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1205: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1206: out = 32'b11010010100111010001110100000001; // MOVZ X1, 59624
         16'd1207: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1208: out = 32'b11110010100100101000101000000001; // MOVK X1, 37968
         16'd1209: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1210: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd1211: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1212: out = 32'b11110010100010101001010100000001; // MOVK X1, 21672
         16'd1213: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1214: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1215: out = 32'b11010010100111010000100000000001; // MOVZ X1, 59456
         16'd1216: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1217: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1218: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1219: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1220: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1221: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1222: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1223: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1224: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1225: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1226: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1227: out = 32'b11010010100000010000000100000001; // MOVZ X1, 2056
         16'd1228: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1229: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd1230: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1231: out = 32'b11110010100000010000000010000001; // MOVK X1, 2052
         16'd1232: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1233: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1234: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1235: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1236: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd1237: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1238: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1239: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1240: out = 32'b11110010100010110000101100000001; // MOVK X1, 22616
         16'd1241: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1242: out = 32'b11110010100000010000001100000001; // MOVK X1, 2072
         16'd1243: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1244: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1245: out = 32'b11010010100000110000101100000001; // MOVZ X1, 6232
         16'd1246: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1247: out = 32'b11110010100010110000001100000001; // MOVK X1, 22552
         16'd1248: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1249: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1250: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1251: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1252: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1253: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1254: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd1255: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1256: out = 32'b11110010100000000000100000000001; // MOVK X1, 64
         16'd1257: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1258: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd1259: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1260: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd1261: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1262: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1263: out = 32'b11010010100100101001001010000001; // MOVZ X1, 38036
         16'd1264: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1265: out = 32'b11110010100101001001110100000001; // MOVK X1, 42216
         16'd1266: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1267: out = 32'b11110010100111010001111100000001; // MOVK X1, 59640
         16'd1268: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1269: out = 32'b11110010100111111001111110000001; // MOVK X1, 64764
         16'd1270: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1271: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1272: out = 32'b11010010100111111001111110000001; // MOVZ X1, 64764
         16'd1273: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1274: out = 32'b11110010100111111001111110000001; // MOVK X1, 64764
         16'd1275: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1276: out = 32'b11110010100111110001111100000001; // MOVK X1, 63736
         16'd1277: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1278: out = 32'b11110010100111110001110100000001; // MOVK X1, 63720
         16'd1279: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1280: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1281: out = 32'b11010010100111010001110100000001; // MOVZ X1, 59624
         16'd1282: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1283: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd1284: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1285: out = 32'b11110010100010101000101010000001; // MOVK X1, 21588
         16'd1286: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1287: out = 32'b11110010100010101001110100000001; // MOVK X1, 21736
         16'd1288: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1289: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1290: out = 32'b11010010100111010000101000000001; // MOVZ X1, 59472
         16'd1291: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1292: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1293: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1294: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1295: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1296: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1297: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1298: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1299: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd1300: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1301: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1302: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1303: out = 32'b11010010100010110000101100000001; // MOVZ X1, 22616
         16'd1304: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1305: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd1306: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1307: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd1308: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1309: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1310: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1311: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1312: out = 32'b11010010100000001000001100000001; // MOVZ X1, 1048
         16'd1313: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1314: out = 32'b11110010100010110000101010000001; // MOVK X1, 22612
         16'd1315: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1316: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1317: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1318: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1319: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1320: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1321: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd1322: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1323: out = 32'b11110010100010000000101010000001; // MOVK X1, 16468
         16'd1324: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1325: out = 32'b11110010100010100000101000000001; // MOVK X1, 20560
         16'd1326: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1327: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd1328: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1329: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1330: out = 32'b11010010100010100000101000000001; // MOVZ X1, 20560
         16'd1331: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1332: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd1333: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1334: out = 32'b11110010100111010001111100000001; // MOVK X1, 59640
         16'd1335: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1336: out = 32'b11110010100111110001111110000001; // MOVK X1, 63740
         16'd1337: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1338: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1339: out = 32'b11010010100111111001111100000001; // MOVZ X1, 64760
         16'd1340: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1341: out = 32'b11110010100111111001111110000001; // MOVK X1, 64764
         16'd1342: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1343: out = 32'b11110010100111110001111100000001; // MOVK X1, 63736
         16'd1344: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1345: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd1346: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1347: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1348: out = 32'b11010010100111010001110100000001; // MOVZ X1, 59624
         16'd1349: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1350: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd1351: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1352: out = 32'b11110010100010101000101010000001; // MOVK X1, 21588
         16'd1353: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1354: out = 32'b11110010100100101001110010000001; // MOVK X1, 38116
         16'd1355: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1356: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1357: out = 32'b11010010100111001001001000000001; // MOVZ X1, 58512
         16'd1358: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1359: out = 32'b11110010100010000000000000000001; // MOVK X1, 16384
         16'd1360: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1361: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1362: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1363: out = 32'b11110010100000000000100000000001; // MOVK X1, 64
         16'd1364: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1365: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1366: out = 32'b11111000000000000000000001001010; // STUR X10, [X2, 0]
         16'd1367: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1368: out = 32'b11010010100000010000000100000001; // MOVZ X1, 2056
         16'd1369: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1370: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd1371: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1372: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd1373: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1374: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1375: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1376: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1377: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd1378: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1379: out = 32'b11110010100010110000101100000001; // MOVK X1, 22616
         16'd1380: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1381: out = 32'b11110010100010010000000100000001; // MOVK X1, 18440
         16'd1382: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1383: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd1384: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1385: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1386: out = 32'b11010010100010110000000100000001; // MOVZ X1, 22536
         16'd1387: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1388: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd1389: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1390: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1391: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1392: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1393: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1394: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1395: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd1396: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1397: out = 32'b11110010100010001000100010000001; // MOVK X1, 17476
         16'd1398: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1399: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1400: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1401: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1402: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1403: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1404: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd1405: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1406: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd1407: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1408: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd1409: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1410: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd1411: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1412: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1413: out = 32'b11010010100010000000100000000001; // MOVZ X1, 16448
         16'd1414: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1415: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd1416: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1417: out = 32'b11110010100100101001110100000001; // MOVK X1, 38120
         16'd1418: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1419: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd1420: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1421: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1422: out = 32'b11010010100111110001111100000001; // MOVZ X1, 63736
         16'd1423: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1424: out = 32'b11110010100111110001111100000001; // MOVK X1, 63736
         16'd1425: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1426: out = 32'b11110010100111110001111100000001; // MOVK X1, 63736
         16'd1427: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1428: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd1429: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1430: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1431: out = 32'b11010010100111010001110100000001; // MOVZ X1, 59624
         16'd1432: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1433: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd1434: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1435: out = 32'b11110010100010101000101000000001; // MOVK X1, 21584
         16'd1436: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1437: out = 32'b11110010100010101001001010000001; // MOVK X1, 21652
         16'd1438: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1439: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1440: out = 32'b11010010100100101001101010000001; // MOVZ X1, 38100
         16'd1441: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1442: out = 32'b11110010100110101000101000000001; // MOVK X1, 54352
         16'd1443: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1444: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1445: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1446: out = 32'b11110010100000000000101000000001; // MOVK X1, 80
         16'd1447: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1448: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1449: out = 32'b11010010100100101001001010000001; // MOVZ X1, 38036
         16'd1450: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1451: out = 32'b11110010100010100000000000000001; // MOVK X1, 20480
         16'd1452: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1453: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1454: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1455: out = 32'b11110010100010000001001000000001; // MOVK X1, 16528
         16'd1456: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1457: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1458: out = 32'b11010010100000010000000100000001; // MOVZ X1, 2056
         16'd1459: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1460: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd1461: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1462: out = 32'b11110010100000010000000010000001; // MOVK X1, 2052
         16'd1463: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1464: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1465: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1466: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1467: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd1468: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1469: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1470: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1471: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1472: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1473: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd1474: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1475: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1476: out = 32'b11010010100000010000000010000001; // MOVZ X1, 2052
         16'd1477: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1478: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1479: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1480: out = 32'b11110010100010001000100010000001; // MOVK X1, 17476
         16'd1481: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1482: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1483: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1484: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1485: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd1486: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1487: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1488: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1489: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd1490: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1491: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1492: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1493: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1494: out = 32'b11010010100000000000101010000001; // MOVZ X1, 84
         16'd1495: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1496: out = 32'b11110010100010101000100000000001; // MOVK X1, 21568
         16'd1497: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1498: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd1499: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1500: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd1501: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1502: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1503: out = 32'b11010010100010000000100000000001; // MOVZ X1, 16448
         16'd1504: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1505: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd1506: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1507: out = 32'b11110010100010000000101000000001; // MOVK X1, 16464
         16'd1508: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1509: out = 32'b11110010100100101001110100000001; // MOVK X1, 38120
         16'd1510: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1511: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1512: out = 32'b11111000000000000000000001010001; // STUR X17, [X2, 0]
         16'd1513: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1514: out = 32'b11010010100111010001110100000001; // MOVZ X1, 59624
         16'd1515: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1516: out = 32'b11110010100100101000101000000001; // MOVK X1, 37968
         16'd1517: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1518: out = 32'b11110010100010000000000000000001; // MOVK X1, 16384
         16'd1519: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1520: out = 32'b11110010100010100001010010000001; // MOVK X1, 20644
         16'd1521: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1522: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1523: out = 32'b11010010100101000001110010000001; // MOVZ X1, 41188
         16'd1524: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1525: out = 32'b11110010100111001001010010000001; // MOVK X1, 58532
         16'd1526: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1527: out = 32'b11110010100011001000110010000001; // MOVK X1, 25700
         16'd1528: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1529: out = 32'b11110010100011001001010010000001; // MOVK X1, 25764
         16'd1530: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1531: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1532: out = 32'b11010010100111001001110010000001; // MOVZ X1, 58596
         16'd1533: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1534: out = 32'b11110010100101001000101000000001; // MOVK X1, 42064
         16'd1535: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1536: out = 32'b11110010100011000000101000000001; // MOVK X1, 24656
         16'd1537: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1538: out = 32'b11110010100100101001110010000001; // MOVK X1, 38116
         16'd1539: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1540: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1541: out = 32'b11010010100000010000000100000001; // MOVZ X1, 2056
         16'd1542: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1543: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd1544: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1545: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1546: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1547: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1548: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1549: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1550: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd1551: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1552: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd1553: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1554: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1555: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1556: out = 32'b11110010100010110000101100000001; // MOVK X1, 22616
         16'd1557: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1558: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1559: out = 32'b11010010100010110000101100000001; // MOVZ X1, 22616
         16'd1560: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1561: out = 32'b11110010100010110000100010000001; // MOVK X1, 22596
         16'd1562: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1563: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1564: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1565: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1566: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1567: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1568: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd1569: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1570: out = 32'b11110010100000001000100010000001; // MOVK X1, 1092
         16'd1571: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1572: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd1573: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1574: out = 32'b11110010100010000000000000000001; // MOVK X1, 16384
         16'd1575: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1576: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1577: out = 32'b11010010100010000001001010000001; // MOVZ X1, 16532
         16'd1578: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1579: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd1580: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1581: out = 32'b11110010100010100000100000000001; // MOVK X1, 20544
         16'd1582: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1583: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd1584: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1585: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1586: out = 32'b11010010100010000000100000000001; // MOVZ X1, 16448
         16'd1587: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1588: out = 32'b11110010100010100000100000000001; // MOVK X1, 20544
         16'd1589: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1590: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd1591: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1592: out = 32'b11110010100100101001110100000001; // MOVK X1, 38120
         16'd1593: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1594: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1595: out = 32'b11010010100111010001110100000001; // MOVZ X1, 59624
         16'd1596: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1597: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd1598: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1599: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd1600: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1601: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd1602: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1603: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1604: out = 32'b11010010100111010001110100000001; // MOVZ X1, 59624
         16'd1605: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1606: out = 32'b11110010100100101000100000000001; // MOVK X1, 37952
         16'd1607: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1608: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1609: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1610: out = 32'b11110010100010100000110010000001; // MOVK X1, 20580
         16'd1611: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1612: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1613: out = 32'b11010010100101001001110010000001; // MOVZ X1, 42212
         16'd1614: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1615: out = 32'b11110010100101001001010010000001; // MOVK X1, 42148
         16'd1616: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1617: out = 32'b11110010100011000000110000000001; // MOVK X1, 24672
         16'd1618: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1619: out = 32'b11110010100011001001010010000001; // MOVK X1, 25764
         16'd1620: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1621: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1622: out = 32'b11010010100111001001110010000001; // MOVZ X1, 58596
         16'd1623: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1624: out = 32'b11110010100111001001010010000001; // MOVK X1, 58532
         16'd1625: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1626: out = 32'b11110010100101101001010010000001; // MOVK X1, 46244
         16'd1627: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1628: out = 32'b11110010100111001001110010000001; // MOVK X1, 58596
         16'd1629: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1630: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1631: out = 32'b11010010100000010000000100000001; // MOVZ X1, 2056
         16'd1632: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1633: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd1634: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1635: out = 32'b11110010100000010000000010000001; // MOVK X1, 2052
         16'd1636: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1637: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1638: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1639: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1640: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd1641: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1642: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1643: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1644: out = 32'b11110010100010101000101100000001; // MOVK X1, 21592
         16'd1645: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1646: out = 32'b11110010100010110000101100000001; // MOVK X1, 22616
         16'd1647: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1648: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1649: out = 32'b11010010100010110000000010000001; // MOVZ X1, 22532
         16'd1650: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1651: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd1652: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1653: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1654: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1655: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1656: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1657: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1658: out = 32'b11010010100000001000101010000001; // MOVZ X1, 1108
         16'd1659: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1660: out = 32'b11110010100010101000100010000001; // MOVK X1, 21572
         16'd1661: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1662: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd1663: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1664: out = 32'b11110010100100101000100000000001; // MOVK X1, 37952
         16'd1665: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1666: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1667: out = 32'b11010010100010000001001010000001; // MOVZ X1, 16532
         16'd1668: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1669: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd1670: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1671: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd1672: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1673: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd1674: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1675: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1676: out = 32'b11010010100100101001110100000001; // MOVZ X1, 38120
         16'd1677: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1678: out = 32'b11110010100111010001010100000001; // MOVK X1, 59560
         16'd1679: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1680: out = 32'b11110010100100101000101000000001; // MOVK X1, 37968
         16'd1681: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1682: out = 32'b11110010100100100001110100000001; // MOVK X1, 37096
         16'd1683: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1684: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1685: out = 32'b11010010100111010001110010000001; // MOVZ X1, 59620
         16'd1686: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1687: out = 32'b11110010100010100000100000000001; // MOVK X1, 20544
         16'd1688: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1689: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd1690: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1691: out = 32'b11110010100100101001010010000001; // MOVK X1, 38052
         16'd1692: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1693: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1694: out = 32'b11010010100111010001110100000001; // MOVZ X1, 59624
         16'd1695: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1696: out = 32'b11110010100010100000000000000001; // MOVK X1, 20480
         16'd1697: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1698: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1699: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1700: out = 32'b11110010100010100000110010000001; // MOVK X1, 20580
         16'd1701: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1702: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1703: out = 32'b11010010100101001001010010000001; // MOVZ X1, 42148
         16'd1704: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1705: out = 32'b11110010100101001001010010000001; // MOVK X1, 42148
         16'd1706: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1707: out = 32'b11110010100011000000110010000001; // MOVK X1, 24676
         16'd1708: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1709: out = 32'b11110010100011001001010010000001; // MOVK X1, 25764
         16'd1710: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1711: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1712: out = 32'b11010010100100100001001000000001; // MOVZ X1, 37008
         16'd1713: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1714: out = 32'b11110010100101001001010010000001; // MOVK X1, 42148
         16'd1715: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1716: out = 32'b11110010100011001001010010000001; // MOVK X1, 25764
         16'd1717: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1718: out = 32'b11110010100101001001010010000001; // MOVK X1, 42148
         16'd1719: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1720: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1721: out = 32'b11010010100000010000000100000001; // MOVZ X1, 2056
         16'd1722: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1723: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd1724: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1725: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd1726: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1727: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1728: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1729: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1730: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd1731: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1732: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1733: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1734: out = 32'b11110010100010110000100010000001; // MOVK X1, 22596
         16'd1735: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1736: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1737: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1738: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1739: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd1740: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1741: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd1742: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1743: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1744: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1745: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd1746: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1747: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1748: out = 32'b11010010100000000000000010000001; // MOVZ X1, 4
         16'd1749: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1750: out = 32'b11110010100000001000100000000001; // MOVK X1, 1088
         16'd1751: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1752: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd1753: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1754: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd1755: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1756: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1757: out = 32'b11010010100100101001001010000001; // MOVZ X1, 38036
         16'd1758: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1759: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd1760: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1761: out = 32'b11110010100100101001010010000001; // MOVK X1, 38052
         16'd1762: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1763: out = 32'b11110010100111001001101010000001; // MOVK X1, 58580
         16'd1764: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1765: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1766: out = 32'b11010010100100101001110010000001; // MOVZ X1, 38116
         16'd1767: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1768: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd1769: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1770: out = 32'b11110010100101001001001010000001; // MOVK X1, 42132
         16'd1771: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1772: out = 32'b11110010100100100001110010000001; // MOVK X1, 37092
         16'd1773: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1774: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1775: out = 32'b11010010100111001001010010000001; // MOVZ X1, 58532
         16'd1776: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1777: out = 32'b11110010100100101000100000000001; // MOVK X1, 37952
         16'd1778: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1779: out = 32'b11110010100010000000101000000001; // MOVK X1, 16464
         16'd1780: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1781: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd1782: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1783: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1784: out = 32'b11010010100111001001010010000001; // MOVZ X1, 58532
         16'd1785: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1786: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1787: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1788: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1789: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1790: out = 32'b11110010100000100000110010000001; // MOVK X1, 4196
         16'd1791: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1792: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1793: out = 32'b11010010100011001000110010000001; // MOVZ X1, 25700
         16'd1794: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1795: out = 32'b11110010100011001000110000000001; // MOVK X1, 25696
         16'd1796: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1797: out = 32'b11110010100011000000110010000001; // MOVK X1, 24676
         16'd1798: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1799: out = 32'b11110010100011001000110010000001; // MOVK X1, 25700
         16'd1800: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1801: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1802: out = 32'b11010010100010100000101000000001; // MOVZ X1, 20560
         16'd1803: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1804: out = 32'b11110010100101001000110010000001; // MOVK X1, 42084
         16'd1805: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1806: out = 32'b11110010100011001000110010000001; // MOVK X1, 25700
         16'd1807: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1808: out = 32'b11110010100011001000110010000001; // MOVK X1, 25700
         16'd1809: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1810: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1811: out = 32'b11010010100000010000000100000001; // MOVZ X1, 2056
         16'd1812: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1813: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd1814: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1815: out = 32'b11110010100000010000000010000001; // MOVK X1, 2052
         16'd1816: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1817: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1818: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1819: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1820: out = 32'b11010010100000001000000000000001; // MOVZ X1, 1024
         16'd1821: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1822: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1823: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1824: out = 32'b11110010100010110000101010000001; // MOVK X1, 22612
         16'd1825: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1826: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1827: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1828: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1829: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd1830: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1831: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1832: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1833: out = 32'b11110010100000001000101010000001; // MOVK X1, 1108
         16'd1834: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1835: out = 32'b11110010100010101000100010000001; // MOVK X1, 21572
         16'd1836: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1837: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1838: out = 32'b11010010100000001000000000000001; // MOVZ X1, 1024
         16'd1839: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1840: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1841: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1842: out = 32'b11110010100100101001001000000001; // MOVK X1, 38032
         16'd1843: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1844: out = 32'b11110010100010000001001000000001; // MOVK X1, 16528
         16'd1845: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1846: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1847: out = 32'b11010010100100101001001010000001; // MOVZ X1, 38036
         16'd1848: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1849: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd1850: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1851: out = 32'b11110010100100101001110010000001; // MOVK X1, 38116
         16'd1852: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1853: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd1854: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1855: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1856: out = 32'b11010010100111010001110100000001; // MOVZ X1, 59624
         16'd1857: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1858: out = 32'b11110010100111010001110010000001; // MOVK X1, 59620
         16'd1859: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1860: out = 32'b11110010100100101001001000000001; // MOVK X1, 38032
         16'd1861: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1862: out = 32'b11110010100100101001110100000001; // MOVK X1, 38120
         16'd1863: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1864: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1865: out = 32'b11010010100111010001010010000001; // MOVZ X1, 59556
         16'd1866: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1867: out = 32'b11110010100111010001010010000001; // MOVK X1, 59556
         16'd1868: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1869: out = 32'b11110010100100101000101000000001; // MOVK X1, 37968
         16'd1870: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1871: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd1872: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1873: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1874: out = 32'b11010010100100101000101010000001; // MOVZ X1, 37972
         16'd1875: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1876: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1877: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1878: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1879: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1880: out = 32'b11110010100000100000110010000001; // MOVK X1, 4196
         16'd1881: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1882: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1883: out = 32'b11111000000000000000000001001111; // STUR X15, [X2, 0]
         16'd1884: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1885: out = 32'b11010010100010100000101000000001; // MOVZ X1, 20560
         16'd1886: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1887: out = 32'b11110010100011001000110010000001; // MOVK X1, 25700
         16'd1888: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1889: out = 32'b11110010100011001000110010000001; // MOVK X1, 25700
         16'd1890: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1891: out = 32'b11110010100011001000110010000001; // MOVK X1, 25700
         16'd1892: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1893: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1894: out = 32'b11010010100000010000000100000001; // MOVZ X1, 2056
         16'd1895: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1896: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd1897: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1898: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1899: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1900: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1901: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1902: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1903: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd1904: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1905: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1906: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1907: out = 32'b11110010100010110000101100000001; // MOVK X1, 22616
         16'd1908: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1909: out = 32'b11110010100010101000000010000001; // MOVK X1, 21508
         16'd1910: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1911: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1912: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd1913: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1914: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1915: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1916: out = 32'b11110010100000001000101010000001; // MOVK X1, 1108
         16'd1917: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1918: out = 32'b11110010100010101000100010000001; // MOVK X1, 21572
         16'd1919: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1920: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1921: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd1922: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1923: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1924: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1925: out = 32'b11110010100100101001001000000001; // MOVK X1, 38032
         16'd1926: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1927: out = 32'b11110010100100100001001010000001; // MOVK X1, 37012
         16'd1928: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1929: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1930: out = 32'b11010010100100100001001010000001; // MOVZ X1, 37012
         16'd1931: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1932: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd1933: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1934: out = 32'b11110010100100101001101010000001; // MOVK X1, 38100
         16'd1935: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1936: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd1937: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1938: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1939: out = 32'b11010010100111010001110100000001; // MOVZ X1, 59624
         16'd1940: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1941: out = 32'b11110010100111001001110010000001; // MOVK X1, 58596
         16'd1942: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1943: out = 32'b11110010100110101001001010000001; // MOVK X1, 54420
         16'd1944: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1945: out = 32'b11110010100111001001110100000001; // MOVK X1, 58600
         16'd1946: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1947: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1948: out = 32'b11010010100111010001110100000001; // MOVZ X1, 59624
         16'd1949: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1950: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd1951: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1952: out = 32'b11110010100111010001010010000001; // MOVK X1, 59556
         16'd1953: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1954: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd1955: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1956: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1957: out = 32'b11010010100100101000100000000001; // MOVZ X1, 37952
         16'd1958: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1959: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1960: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1961: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd1962: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1963: out = 32'b11110010100010100000110010000001; // MOVK X1, 20580
         16'd1964: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1965: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1966: out = 32'b11010010100101000001010000000001; // MOVZ X1, 41120
         16'd1967: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1968: out = 32'b11110010100101000000110000000001; // MOVK X1, 41056
         16'd1969: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1970: out = 32'b11110010100011001000110010000001; // MOVK X1, 25700
         16'd1971: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1972: out = 32'b11110010100011001001010010000001; // MOVK X1, 25764
         16'd1973: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1974: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1975: out = 32'b11010010100010100000100000000001; // MOVZ X1, 20544
         16'd1976: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1977: out = 32'b11110010100000100000001000000001; // MOVK X1, 4112
         16'd1978: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1979: out = 32'b11110010100010100000110010000001; // MOVK X1, 20580
         16'd1980: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1981: out = 32'b11110010100011000000101000000001; // MOVK X1, 24656
         16'd1982: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1983: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1984: out = 32'b11010010100000010000000100000001; // MOVZ X1, 2056
         16'd1985: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1986: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd1987: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1988: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd1989: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1990: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1991: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd1992: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd1993: out = 32'b11010010100000000000000010000001; // MOVZ X1, 4
         16'd1994: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1995: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd1996: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1997: out = 32'b11110010100010110000101100000001; // MOVK X1, 22616
         16'd1998: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd1999: out = 32'b11110010100010101000000010000001; // MOVK X1, 21508
         16'd2000: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2001: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2002: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd2003: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2004: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd2005: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2006: out = 32'b11110010100000001000101010000001; // MOVK X1, 1108
         16'd2007: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2008: out = 32'b11110010100010101000101010000001; // MOVK X1, 21588
         16'd2009: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2010: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2011: out = 32'b11010010100010001000000010000001; // MOVZ X1, 17412
         16'd2012: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2013: out = 32'b11110010100010101000100000000001; // MOVK X1, 21568
         16'd2014: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2015: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd2016: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2017: out = 32'b11110010100100101001001000000001; // MOVK X1, 38032
         16'd2018: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2019: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2020: out = 32'b11010010100100100001001000000001; // MOVZ X1, 37008
         16'd2021: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2022: out = 32'b11110010100100100001001000000001; // MOVK X1, 37008
         16'd2023: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2024: out = 32'b11110010100100101001101010000001; // MOVK X1, 38100
         16'd2025: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2026: out = 32'b11110010100111001001110100000001; // MOVK X1, 58600
         16'd2027: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2028: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2029: out = 32'b11010010100111010001001010000001; // MOVZ X1, 59540
         16'd2030: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2031: out = 32'b11110010100100101001101010000001; // MOVK X1, 38100
         16'd2032: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2033: out = 32'b11110010100110101001101010000001; // MOVK X1, 54484
         16'd2034: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2035: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd2036: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2037: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2038: out = 32'b11010010100111110001110100000001; // MOVZ X1, 63720
         16'd2039: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2040: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd2041: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2042: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd2043: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2044: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd2045: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2046: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2047: out = 32'b11010010100010101000000000000001; // MOVZ X1, 21504
         16'd2048: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2049: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2050: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2051: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2052: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2053: out = 32'b11110010100011001001010000000001; // MOVK X1, 25760
         16'd2054: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2055: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2056: out = 32'b11010010100101100001110000000001; // MOVZ X1, 45280
         16'd2057: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2058: out = 32'b11110010100111000001011000000001; // MOVK X1, 57520
         16'd2059: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2060: out = 32'b11110010100011000000110010000001; // MOVK X1, 24676
         16'd2061: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2062: out = 32'b11110010100011000001010010000001; // MOVK X1, 24740
         16'd2063: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2064: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2065: out = 32'b11010010100101000001001010000001; // MOVZ X1, 41108
         16'd2066: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2067: out = 32'b11110010100010000000000000000001; // MOVK X1, 16384
         16'd2068: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2069: out = 32'b11110010100000100001011100000001; // MOVK X1, 4280
         16'd2070: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2071: out = 32'b11110010100101001001001000000001; // MOVK X1, 42128
         16'd2072: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2073: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2074: out = 32'b11010010100000010000000100000001; // MOVZ X1, 2056
         16'd2075: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2076: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd2077: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2078: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd2079: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2080: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd2081: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2082: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2083: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd2084: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2085: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd2086: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2087: out = 32'b11110010100010110000101010000001; // MOVK X1, 22612
         16'd2088: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2089: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd2090: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2091: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2092: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd2093: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2094: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd2095: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2096: out = 32'b11110010100000001000101010000001; // MOVK X1, 1108
         16'd2097: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2098: out = 32'b11110010100010110000101010000001; // MOVK X1, 22612
         16'd2099: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2100: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2101: out = 32'b11010010100010001000000010000001; // MOVZ X1, 17412
         16'd2102: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2103: out = 32'b11110010100010101000100000000001; // MOVK X1, 21568
         16'd2104: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2105: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd2106: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2107: out = 32'b11110010100100101001001000000001; // MOVK X1, 38032
         16'd2108: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2109: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2110: out = 32'b11010010100100100001001000000001; // MOVZ X1, 37008
         16'd2111: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2112: out = 32'b11110010100100100001001000000001; // MOVK X1, 37008
         16'd2113: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2114: out = 32'b11110010100100101001101010000001; // MOVK X1, 38100
         16'd2115: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2116: out = 32'b11110010100111001001110100000001; // MOVK X1, 58600
         16'd2117: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2118: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2119: out = 32'b11010010100100101000100000000001; // MOVZ X1, 37952
         16'd2120: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2121: out = 32'b11110010100100101001110010000001; // MOVK X1, 38116
         16'd2122: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2123: out = 32'b11110010100111001001101010000001; // MOVK X1, 58580
         16'd2124: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2125: out = 32'b11110010100111010001111100000001; // MOVK X1, 59640
         16'd2126: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2127: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2128: out = 32'b11010010100111110001110100000001; // MOVZ X1, 63720
         16'd2129: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2130: out = 32'b11110010100111010001111100000001; // MOVK X1, 59640
         16'd2131: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2132: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd2133: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2134: out = 32'b11110010100111010001001010000001; // MOVK X1, 59540
         16'd2135: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2136: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2137: out = 32'b11010010100010101000000000000001; // MOVZ X1, 21504
         16'd2138: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2139: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2140: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2141: out = 32'b11110010100000000000001000000001; // MOVK X1, 16
         16'd2142: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2143: out = 32'b11110010100011001001010010000001; // MOVK X1, 25764
         16'd2144: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2145: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2146: out = 32'b11010010100111000001110000000001; // MOVZ X1, 57568
         16'd2147: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2148: out = 32'b11110010100111000001010000000001; // MOVK X1, 57504
         16'd2149: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2150: out = 32'b11110010100011000000110010000001; // MOVK X1, 24676
         16'd2151: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2152: out = 32'b11110010100011000001010000000001; // MOVK X1, 24736
         16'd2153: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2154: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2155: out = 32'b11010010100111001001110010000001; // MOVZ X1, 58596
         16'd2156: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2157: out = 32'b11110010100100100000000000000001; // MOVK X1, 36864
         16'd2158: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2159: out = 32'b11110010100011001001010010000001; // MOVK X1, 25764
         16'd2160: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2161: out = 32'b11110010100111001001110010000001; // MOVK X1, 58596
         16'd2162: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2163: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2164: out = 32'b11010010100000001000000100000001; // MOVZ X1, 1032
         16'd2165: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2166: out = 32'b11110010100000010000000100000001; // MOVK X1, 2056
         16'd2167: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2168: out = 32'b11110010100000010000000010000001; // MOVK X1, 2052
         16'd2169: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2170: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd2171: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2172: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2173: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd2174: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2175: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd2176: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2177: out = 32'b11110010100010110000101100000001; // MOVK X1, 22616
         16'd2178: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2179: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd2180: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2181: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2182: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd2183: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2184: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2185: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2186: out = 32'b11110010100000001000101010000001; // MOVK X1, 1108
         16'd2187: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2188: out = 32'b11110010100010110000101010000001; // MOVK X1, 22612
         16'd2189: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2190: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2191: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd2192: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2193: out = 32'b11110010100010001000100000000001; // MOVK X1, 17472
         16'd2194: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2195: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd2196: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2197: out = 32'b11110010100100101000101000000001; // MOVK X1, 37968
         16'd2198: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2199: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2200: out = 32'b11010010100010100001001000000001; // MOVZ X1, 20624
         16'd2201: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2202: out = 32'b11110010100100100001001000000001; // MOVK X1, 37008
         16'd2203: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2204: out = 32'b11110010100100101001101010000001; // MOVK X1, 38100
         16'd2205: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2206: out = 32'b11110010100111001001110010000001; // MOVK X1, 58596
         16'd2207: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2208: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2209: out = 32'b11010010100100100000100000000001; // MOVZ X1, 36928
         16'd2210: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2211: out = 32'b11110010100010000001001010000001; // MOVK X1, 16532
         16'd2212: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2213: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd2214: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2215: out = 32'b11110010100111010001111100000001; // MOVK X1, 59640
         16'd2216: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2217: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2218: out = 32'b11010010100111110001110100000001; // MOVZ X1, 63720
         16'd2219: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2220: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd2221: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2222: out = 32'b11110010100111110001111100000001; // MOVK X1, 63736
         16'd2223: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2224: out = 32'b11110010100111010001010010000001; // MOVK X1, 59556
         16'd2225: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2226: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2227: out = 32'b11010010100101001000100000000001; // MOVZ X1, 42048
         16'd2228: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2229: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2230: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2231: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2232: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2233: out = 32'b11110010100011001001010010000001; // MOVK X1, 25764
         16'd2234: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2235: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2236: out = 32'b11010010100101000001110000000001; // MOVZ X1, 41184
         16'd2237: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2238: out = 32'b11110010100111000001010000000001; // MOVK X1, 57504
         16'd2239: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2240: out = 32'b11110010100011001000110010000001; // MOVK X1, 25700
         16'd2241: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2242: out = 32'b11110010100011001001010010000001; // MOVK X1, 25764
         16'd2243: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2244: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2245: out = 32'b11010010100111001001110010000001; // MOVZ X1, 58596
         16'd2246: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2247: out = 32'b11110010100100100000101000000001; // MOVK X1, 36944
         16'd2248: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2249: out = 32'b11110010100011001001011100000001; // MOVK X1, 25784
         16'd2250: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2251: out = 32'b11110010100111001001110010000001; // MOVK X1, 58596
         16'd2252: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2253: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2254: out = 32'b11111000000000000000000001010011; // STUR X19, [X2, 0]
         16'd2255: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2256: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd2257: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2258: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd2259: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2260: out = 32'b11110010100010110000101100000001; // MOVK X1, 22616
         16'd2261: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2262: out = 32'b11110010100010110000000010000001; // MOVK X1, 22532
         16'd2263: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2264: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2265: out = 32'b11010010100000001000000000000001; // MOVZ X1, 1024
         16'd2266: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2267: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2268: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2269: out = 32'b11110010100000000000101010000001; // MOVK X1, 84
         16'd2270: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2271: out = 32'b11110010100010101000000000000001; // MOVK X1, 21504
         16'd2272: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2273: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2274: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd2275: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2276: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2277: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2278: out = 32'b11110010100010000000101000000001; // MOVK X1, 16464
         16'd2279: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2280: out = 32'b11110010100010100000101000000001; // MOVK X1, 20560
         16'd2281: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2282: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2283: out = 32'b11010010100010100000101000000001; // MOVZ X1, 20560
         16'd2284: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2285: out = 32'b11110010100010100001001000000001; // MOVK X1, 20624
         16'd2286: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2287: out = 32'b11110010100100101001110010000001; // MOVK X1, 38116
         16'd2288: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2289: out = 32'b11110010100111001001001010000001; // MOVK X1, 58516
         16'd2290: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2291: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2292: out = 32'b11010010100010000000100000000001; // MOVZ X1, 16448
         16'd2293: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2294: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2295: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2296: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd2297: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2298: out = 32'b11110010100100101001110100000001; // MOVK X1, 38120
         16'd2299: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2300: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2301: out = 32'b11010010100111010001110100000001; // MOVZ X1, 59624
         16'd2302: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2303: out = 32'b11110010100111001001001010000001; // MOVK X1, 58516
         16'd2304: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2305: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd2306: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2307: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd2308: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2309: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2310: out = 32'b11010010100101010000000000000001; // MOVZ X1, 43008
         16'd2311: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2312: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2313: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2314: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2315: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2316: out = 32'b11110010100000100000110010000001; // MOVK X1, 4196
         16'd2317: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2318: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2319: out = 32'b11010010100101001001010000000001; // MOVZ X1, 42144
         16'd2320: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2321: out = 32'b11110010100101001001010010000001; // MOVK X1, 42148
         16'd2322: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2323: out = 32'b11110010100011001000110010000001; // MOVK X1, 25700
         16'd2324: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2325: out = 32'b11110010100011001001010010000001; // MOVK X1, 25764
         16'd2326: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2327: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2328: out = 32'b11010010100100100001001000000001; // MOVZ X1, 37008
         16'd2329: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2330: out = 32'b11110010100101001000001000000001; // MOVK X1, 42000
         16'd2331: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2332: out = 32'b11110010100010101001111100000001; // MOVK X1, 21752
         16'd2333: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2334: out = 32'b11110010100111001001110010000001; // MOVK X1, 58596
         16'd2335: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2336: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2337: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd2338: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2339: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd2340: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2341: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd2342: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2343: out = 32'b11110010100010110000101100000001; // MOVK X1, 22616
         16'd2344: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2345: out = 32'b11110010100010110000000000000001; // MOVK X1, 22528
         16'd2346: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2347: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2348: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd2349: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2350: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2351: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2352: out = 32'b11110010100000000000000010000001; // MOVK X1, 4
         16'd2353: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2354: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2355: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2356: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2357: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd2358: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2359: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2360: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2361: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2362: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2363: out = 32'b11110010100010100000101000000001; // MOVK X1, 20560
         16'd2364: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2365: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2366: out = 32'b11010010100010100000100000000001; // MOVZ X1, 20544
         16'd2367: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2368: out = 32'b11110010100010000001001000000001; // MOVK X1, 16528
         16'd2369: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2370: out = 32'b11110010100100101001101010000001; // MOVK X1, 38100
         16'd2371: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2372: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd2373: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2374: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2375: out = 32'b11010010100010100000100000000001; // MOVZ X1, 20544
         16'd2376: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2377: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2378: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2379: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2380: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2381: out = 32'b11110010100010000001001010000001; // MOVK X1, 16532
         16'd2382: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2383: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2384: out = 32'b11010010100100101001001010000001; // MOVZ X1, 38036
         16'd2385: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2386: out = 32'b11110010100111010001110010000001; // MOVK X1, 59620
         16'd2387: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2388: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd2389: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2390: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd2391: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2392: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2393: out = 32'b11010010100101001000101000000001; // MOVZ X1, 42064
         16'd2394: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2395: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2396: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2397: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2398: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2399: out = 32'b11110010100000100000110010000001; // MOVK X1, 4196
         16'd2400: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2401: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2402: out = 32'b11010010100011001001011010000001; // MOVZ X1, 25780
         16'd2403: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2404: out = 32'b11110010100011000000110000000001; // MOVK X1, 24672
         16'd2405: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2406: out = 32'b11110010100011000000110010000001; // MOVK X1, 24676
         16'd2407: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2408: out = 32'b11110010100011001000110000000001; // MOVK X1, 25696
         16'd2409: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2410: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2411: out = 32'b11010010100011000000101000000001; // MOVZ X1, 24656
         16'd2412: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2413: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2414: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2415: out = 32'b11110010100010101000101010000001; // MOVK X1, 21588
         16'd2416: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2417: out = 32'b11110010100010100001001000000001; // MOVK X1, 20624
         16'd2418: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2419: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2420: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd2421: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2422: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd2423: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2424: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd2425: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2426: out = 32'b11110010100010110000101100000001; // MOVK X1, 22616
         16'd2427: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2428: out = 32'b11110010100010101000000000000001; // MOVK X1, 21504
         16'd2429: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2430: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2431: out = 32'b11010010100000001000000000000001; // MOVZ X1, 1024
         16'd2432: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2433: out = 32'b11110010100000000000000010000001; // MOVK X1, 4
         16'd2434: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2435: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd2436: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2437: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2438: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2439: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2440: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd2441: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2442: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2443: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2444: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2445: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2446: out = 32'b11110010100010100000101000000001; // MOVK X1, 20560
         16'd2447: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2448: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2449: out = 32'b11010010100010100000100000000001; // MOVZ X1, 20544
         16'd2450: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2451: out = 32'b11110010100010000000101000000001; // MOVK X1, 16464
         16'd2452: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2453: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd2454: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2455: out = 32'b11110010100100100000101000000001; // MOVK X1, 36944
         16'd2456: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2457: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2458: out = 32'b11010010100100101001001010000001; // MOVZ X1, 38036
         16'd2459: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2460: out = 32'b11110010100100101000100000000001; // MOVK X1, 37952
         16'd2461: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2462: out = 32'b11110010100010000000101010000001; // MOVK X1, 16468
         16'd2463: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2464: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd2465: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2466: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2467: out = 32'b11010010100101001001110100000001; // MOVZ X1, 42216
         16'd2468: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2469: out = 32'b11110010100111010001110010000001; // MOVK X1, 59620
         16'd2470: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2471: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd2472: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2473: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd2474: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2475: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2476: out = 32'b11010010100111010001001010000001; // MOVZ X1, 59540
         16'd2477: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2478: out = 32'b11110010100000000000100000000001; // MOVK X1, 64
         16'd2479: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2480: out = 32'b11110010100010100000101010000001; // MOVK X1, 20564
         16'd2481: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2482: out = 32'b11110010100010101000110010000001; // MOVK X1, 21604
         16'd2483: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2484: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2485: out = 32'b11010010100101001001010010000001; // MOVZ X1, 42148
         16'd2486: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2487: out = 32'b11110010100011001000110000000001; // MOVK X1, 25696
         16'd2488: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2489: out = 32'b11110010100011000000110010000001; // MOVK X1, 24676
         16'd2490: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2491: out = 32'b11110010100011001000110010000001; // MOVK X1, 25700
         16'd2492: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2493: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2494: out = 32'b11010010100101001000101000000001; // MOVZ X1, 42064
         16'd2495: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2496: out = 32'b11110010100000100000001000000001; // MOVK X1, 4112
         16'd2497: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2498: out = 32'b11110010100101001001111100000001; // MOVK X1, 42232
         16'd2499: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2500: out = 32'b11110010100101001001010010000001; // MOVK X1, 42148
         16'd2501: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2502: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2503: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd2504: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2505: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd2506: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2507: out = 32'b11110010100000000000000010000001; // MOVK X1, 4
         16'd2508: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2509: out = 32'b11110010100010101000101010000001; // MOVK X1, 21588
         16'd2510: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2511: out = 32'b11110010100000000000000010000001; // MOVK X1, 4
         16'd2512: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2513: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2514: out = 32'b11010010100010001000101010000001; // MOVZ X1, 17492
         16'd2515: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2516: out = 32'b11110010100010101000101100000001; // MOVK X1, 21592
         16'd2517: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2518: out = 32'b11110010100010110000101010000001; // MOVK X1, 22612
         16'd2519: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2520: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd2521: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2522: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2523: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd2524: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2525: out = 32'b11110010100010001000000000000001; // MOVK X1, 17408
         16'd2526: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2527: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2528: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2529: out = 32'b11110010100010100000101000000001; // MOVK X1, 20560
         16'd2530: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2531: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2532: out = 32'b11010010100010000000100000000001; // MOVZ X1, 16448
         16'd2533: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2534: out = 32'b11110010100010000000101000000001; // MOVK X1, 16464
         16'd2535: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2536: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd2537: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2538: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd2539: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2540: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2541: out = 32'b11010010100010000000100000000001; // MOVZ X1, 16448
         16'd2542: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2543: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd2544: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2545: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd2546: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2547: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd2548: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2549: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2550: out = 32'b11010010100111010001110100000001; // MOVZ X1, 59624
         16'd2551: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2552: out = 32'b11110010100111010001110010000001; // MOVK X1, 59620
         16'd2553: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2554: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd2555: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2556: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd2557: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2558: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2559: out = 32'b11010010100111010000101010000001; // MOVZ X1, 59476
         16'd2560: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2561: out = 32'b11110010100010000000101000000001; // MOVK X1, 16464
         16'd2562: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2563: out = 32'b11110010100010100000101010000001; // MOVK X1, 20564
         16'd2564: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2565: out = 32'b11110010100011001000101010000001; // MOVK X1, 25684
         16'd2566: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2567: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2568: out = 32'b11010010100101001001010010000001; // MOVZ X1, 42148
         16'd2569: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2570: out = 32'b11110010100010100000101000000001; // MOVK X1, 20560
         16'd2571: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2572: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2573: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2574: out = 32'b11110010100010101000101000000001; // MOVK X1, 21584
         16'd2575: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2576: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2577: out = 32'b11010010100011000000101000000001; // MOVZ X1, 24656
         16'd2578: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2579: out = 32'b11110010100010100000101010000001; // MOVK X1, 20564
         16'd2580: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2581: out = 32'b11110010100011001001010010000001; // MOVK X1, 25764
         16'd2582: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2583: out = 32'b11110010100101001001010010000001; // MOVK X1, 42148
         16'd2584: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2585: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2586: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd2587: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2588: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd2589: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2590: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2591: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2592: out = 32'b11110010100010001000101010000001; // MOVK X1, 17492
         16'd2593: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2594: out = 32'b11110010100000001000101100000001; // MOVK X1, 1112
         16'd2595: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2596: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2597: out = 32'b11010010100010110000101100000001; // MOVZ X1, 22616
         16'd2598: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2599: out = 32'b11110010100010110000101100000001; // MOVK X1, 22616
         16'd2600: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2601: out = 32'b11110010100010110000101100000001; // MOVK X1, 22616
         16'd2602: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2603: out = 32'b11110010100010110000000010000001; // MOVK X1, 22532
         16'd2604: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2605: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2606: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd2607: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2608: out = 32'b11110010100010101000101100000001; // MOVK X1, 21592
         16'd2609: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2610: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2611: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2612: out = 32'b11110010100010000000101000000001; // MOVK X1, 16464
         16'd2613: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2614: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2615: out = 32'b11010010100010000000100000000001; // MOVZ X1, 16448
         16'd2616: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2617: out = 32'b11110010100010000001001000000001; // MOVK X1, 16528
         16'd2618: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2619: out = 32'b11110010100100101001110010000001; // MOVK X1, 38116
         16'd2620: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2621: out = 32'b11110010100010100000100000000001; // MOVK X1, 20544
         16'd2622: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2623: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2624: out = 32'b11010010100010000001001010000001; // MOVZ X1, 16532
         16'd2625: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2626: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd2627: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2628: out = 32'b11110010100100101001101010000001; // MOVK X1, 38100
         16'd2629: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2630: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd2631: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2632: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2633: out = 32'b11010010100111010001110100000001; // MOVZ X1, 59624
         16'd2634: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2635: out = 32'b11110010100111001001110010000001; // MOVK X1, 58596
         16'd2636: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2637: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd2638: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2639: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd2640: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2641: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2642: out = 32'b11010010100111010000100000000001; // MOVZ X1, 59456
         16'd2643: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2644: out = 32'b11110010100100100001110010000001; // MOVK X1, 37092
         16'd2645: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2646: out = 32'b11110010100010100000101010000001; // MOVK X1, 20564
         16'd2647: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2648: out = 32'b11110010100111111001010100000001; // MOVK X1, 64680
         16'd2649: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2650: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2651: out = 32'b11010010100111001001110010000001; // MOVZ X1, 58596
         16'd2652: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2653: out = 32'b11110010100111001001001000000001; // MOVK X1, 58512
         16'd2654: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2655: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd2656: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2657: out = 32'b11110010100010000001001000000001; // MOVK X1, 16528
         16'd2658: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2659: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2660: out = 32'b11010010100110101001001010000001; // MOVZ X1, 54420
         16'd2661: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2662: out = 32'b11110010100010100000000000000001; // MOVK X1, 20480
         16'd2663: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2664: out = 32'b11110010100010100001001010000001; // MOVK X1, 20628
         16'd2665: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2666: out = 32'b11110010100100100001001000000001; // MOVK X1, 37008
         16'd2667: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2668: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2669: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd2670: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2671: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd2672: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2673: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2674: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2675: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd2676: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2677: out = 32'b11110010100000001000101100000001; // MOVK X1, 1112
         16'd2678: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2679: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2680: out = 32'b11010010100010110000101100000001; // MOVZ X1, 22616
         16'd2681: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2682: out = 32'b11110010100010110000101100000001; // MOVK X1, 22616
         16'd2683: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2684: out = 32'b11110010100010110000101100000001; // MOVK X1, 22616
         16'd2685: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2686: out = 32'b11110010100010101000000010000001; // MOVK X1, 21508
         16'd2687: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2688: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2689: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd2690: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2691: out = 32'b11110010100000001001010100000001; // MOVK X1, 1192
         16'd2692: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2693: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2694: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2695: out = 32'b11110010100010100000101000000001; // MOVK X1, 20560
         16'd2696: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2697: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2698: out = 32'b11010010100010000000100000000001; // MOVZ X1, 16448
         16'd2699: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2700: out = 32'b11110010100010000001001000000001; // MOVK X1, 16528
         16'd2701: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2702: out = 32'b11110010100100101001110010000001; // MOVK X1, 38116
         16'd2703: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2704: out = 32'b11110010100110101001001010000001; // MOVK X1, 54420
         16'd2705: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2706: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2707: out = 32'b11010010100100101001001010000001; // MOVZ X1, 38036
         16'd2708: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2709: out = 32'b11110010100101001001110100000001; // MOVK X1, 42216
         16'd2710: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2711: out = 32'b11110010100111111001111110000001; // MOVK X1, 64764
         16'd2712: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2713: out = 32'b11110010100111010001010010000001; // MOVK X1, 59556
         16'd2714: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2715: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2716: out = 32'b11010010100100100001001010000001; // MOVZ X1, 37012
         16'd2717: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2718: out = 32'b11110010100111001001110010000001; // MOVK X1, 58596
         16'd2719: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2720: out = 32'b11110010100111010001110010000001; // MOVK X1, 59620
         16'd2721: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2722: out = 32'b11110010100111001001110100000001; // MOVK X1, 58600
         16'd2723: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2724: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2725: out = 32'b11010010100111010000100000000001; // MOVZ X1, 59456
         16'd2726: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2727: out = 32'b11110010100100101001110010000001; // MOVK X1, 38116
         16'd2728: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2729: out = 32'b11110010100100100000101010000001; // MOVK X1, 36948
         16'd2730: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2731: out = 32'b11110010100101010001010010000001; // MOVK X1, 43172
         16'd2732: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2733: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2734: out = 32'b11010010100111001001110010000001; // MOVZ X1, 58596
         16'd2735: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2736: out = 32'b11110010100111001001001000000001; // MOVK X1, 58512
         16'd2737: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2738: out = 32'b11110010100010101000100000000001; // MOVK X1, 21568
         16'd2739: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2740: out = 32'b11110010100000000001001000000001; // MOVK X1, 144
         16'd2741: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2742: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2743: out = 32'b11010010100111001001110010000001; // MOVZ X1, 58596
         16'd2744: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2745: out = 32'b11110010100101001000000000000001; // MOVK X1, 41984
         16'd2746: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2747: out = 32'b11110010100000000001110100000001; // MOVK X1, 232
         16'd2748: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2749: out = 32'b11110010100111001001110010000001; // MOVK X1, 58596
         16'd2750: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2751: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2752: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd2753: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2754: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd2755: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2756: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2757: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2758: out = 32'b11110010100000000000000010000001; // MOVK X1, 4
         16'd2759: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2760: out = 32'b11110010100000001000101010000001; // MOVK X1, 1108
         16'd2761: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2762: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2763: out = 32'b11010010100010110000101100000001; // MOVZ X1, 22616
         16'd2764: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2765: out = 32'b11110010100010110000101100000001; // MOVK X1, 22616
         16'd2766: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2767: out = 32'b11110010100010110000100010000001; // MOVK X1, 22596
         16'd2768: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2769: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd2770: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2771: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2772: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd2773: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2774: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2775: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2776: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2777: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2778: out = 32'b11110010100010101000100000000001; // MOVK X1, 21568
         16'd2779: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2780: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2781: out = 32'b11010010100010000000100000000001; // MOVZ X1, 16448
         16'd2782: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2783: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd2784: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2785: out = 32'b11110010100100101001101010000001; // MOVK X1, 38100
         16'd2786: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2787: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd2788: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2789: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2790: out = 32'b11010010100100101001001010000001; // MOVZ X1, 38036
         16'd2791: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2792: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd2793: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2794: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd2795: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2796: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd2797: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2798: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2799: out = 32'b11010010100100101001010010000001; // MOVZ X1, 38052
         16'd2800: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2801: out = 32'b11110010100111001001110010000001; // MOVK X1, 58596
         16'd2802: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2803: out = 32'b11110010100111001001110010000001; // MOVK X1, 58596
         16'd2804: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2805: out = 32'b11110010100101001001110100000001; // MOVK X1, 42216
         16'd2806: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2807: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2808: out = 32'b11010010100101001000100000000001; // MOVZ X1, 42048
         16'd2809: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2810: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd2811: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2812: out = 32'b11110010100010000000000000000001; // MOVK X1, 16384
         16'd2813: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2814: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2815: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2816: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2817: out = 32'b11010010100100100001101010000001; // MOVZ X1, 37076
         16'd2818: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2819: out = 32'b11110010100100101000101000000001; // MOVK X1, 37968
         16'd2820: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2821: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2822: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2823: out = 32'b11110010100000000001001000000001; // MOVK X1, 144
         16'd2824: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2825: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2826: out = 32'b11010010100111001001110010000001; // MOVZ X1, 58596
         16'd2827: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2828: out = 32'b11110010100111001000101010000001; // MOVK X1, 58452
         16'd2829: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2830: out = 32'b11110010100000000000101000000001; // MOVK X1, 80
         16'd2831: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2832: out = 32'b11110010100100100001110010000001; // MOVK X1, 37092
         16'd2833: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2834: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2835: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd2836: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2837: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd2838: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2839: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2840: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2841: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2842: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2843: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd2844: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2845: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2846: out = 32'b11010010100010001000101100000001; // MOVZ X1, 17496
         16'd2847: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2848: out = 32'b11110010100010110000101010000001; // MOVK X1, 22612
         16'd2849: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2850: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd2851: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2852: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd2853: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2854: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2855: out = 32'b11010010100000001000000000000001; // MOVZ X1, 1024
         16'd2856: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2857: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2858: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2859: out = 32'b11110010100000000000100000000001; // MOVK X1, 64
         16'd2860: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2861: out = 32'b11110010100100101000100000000001; // MOVK X1, 37952
         16'd2862: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2863: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2864: out = 32'b11010010100010000000100000000001; // MOVZ X1, 16448
         16'd2865: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2866: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd2867: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2868: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd2869: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2870: out = 32'b11110010100100101001001000000001; // MOVK X1, 38032
         16'd2871: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2872: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2873: out = 32'b11010010100100101001101010000001; // MOVZ X1, 38100
         16'd2874: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2875: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd2876: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2877: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd2878: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2879: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd2880: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2881: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2882: out = 32'b11010010100111010001110100000001; // MOVZ X1, 59624
         16'd2883: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2884: out = 32'b11110010100111010001110010000001; // MOVK X1, 59620
         16'd2885: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2886: out = 32'b11110010100111001001010010000001; // MOVK X1, 58532
         16'd2887: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2888: out = 32'b11110010100010101000100000000001; // MOVK X1, 21568
         16'd2889: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2890: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2891: out = 32'b11010010100000000000101000000001; // MOVZ X1, 80
         16'd2892: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2893: out = 32'b11110010100010100000101000000001; // MOVK X1, 20560
         16'd2894: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2895: out = 32'b11110010100010100000001000000001; // MOVK X1, 20496
         16'd2896: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2897: out = 32'b11110010100000100000001000000001; // MOVK X1, 4112
         16'd2898: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2899: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2900: out = 32'b11010010100010100000101000000001; // MOVZ X1, 20560
         16'd2901: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2902: out = 32'b11110010100010100000101000000001; // MOVK X1, 20560
         16'd2903: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2904: out = 32'b11110010100000100000000000000001; // MOVK X1, 4096
         16'd2905: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2906: out = 32'b11110010100010100000101010000001; // MOVK X1, 20564
         16'd2907: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2908: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2909: out = 32'b11010010100111110001110100000001; // MOVZ X1, 63720
         16'd2910: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2911: out = 32'b11110010100111110001010100000001; // MOVK X1, 63656
         16'd2912: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2913: out = 32'b11110010100010101001010100000001; // MOVK X1, 21672
         16'd2914: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2915: out = 32'b11110010100101001001001000000001; // MOVK X1, 42128
         16'd2916: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2917: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2918: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd2919: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2920: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd2921: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2922: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd2923: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2924: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd2925: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2926: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd2927: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2928: out = 32'b11110010100000001000101100000001; // MOVK X1, 1112
         16'd2929: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2930: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2931: out = 32'b11010010100010110000000010000001; // MOVZ X1, 22532
         16'd2932: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2933: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd2934: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2935: out = 32'b11110010100000000000100000000001; // MOVK X1, 64
         16'd2936: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2937: out = 32'b11110010100100101000100000000001; // MOVK X1, 37952
         16'd2938: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2939: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2940: out = 32'b11010010100010000000100000000001; // MOVZ X1, 16448
         16'd2941: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2942: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd2943: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2944: out = 32'b11110010100100100001001010000001; // MOVK X1, 37012
         16'd2945: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2946: out = 32'b11110010100100100001000000000001; // MOVK X1, 36992
         16'd2947: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2948: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2949: out = 32'b11010010100100100001001010000001; // MOVZ X1, 37012
         16'd2950: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2951: out = 32'b11110010100110101001110100000001; // MOVK X1, 54504
         16'd2952: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2953: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd2954: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2955: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd2956: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2957: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2958: out = 32'b11010010100111010001110100000001; // MOVZ X1, 59624
         16'd2959: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2960: out = 32'b11110010100111010001110010000001; // MOVK X1, 59620
         16'd2961: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2962: out = 32'b11110010100101001001001010000001; // MOVK X1, 42132
         16'd2963: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2964: out = 32'b11110010100010000000000000000001; // MOVK X1, 16384
         16'd2965: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2966: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2967: out = 32'b11010010100010100000101000000001; // MOVZ X1, 20560
         16'd2968: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2969: out = 32'b11110010100010101000101000000001; // MOVK X1, 21584
         16'd2970: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2971: out = 32'b11110010100010100000001000000001; // MOVK X1, 20496
         16'd2972: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2973: out = 32'b11110010100000100000001000000001; // MOVK X1, 4112
         16'd2974: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2975: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2976: out = 32'b11010010100010100000101000000001; // MOVZ X1, 20560
         16'd2977: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2978: out = 32'b11110010100010100000001000000001; // MOVK X1, 20496
         16'd2979: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2980: out = 32'b11110010100000100000001000000001; // MOVK X1, 4112
         16'd2981: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2982: out = 32'b11110010100010101000110010000001; // MOVK X1, 21604
         16'd2983: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2984: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2985: out = 32'b11010010100101001001010100000001; // MOVZ X1, 42152
         16'd2986: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2987: out = 32'b11110010100101010000110010000001; // MOVK X1, 43108
         16'd2988: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2989: out = 32'b11110010100011001001011100000001; // MOVK X1, 25784
         16'd2990: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd2991: out = 32'b11110010100101010001001000000001; // MOVK X1, 43152
         16'd2992: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd2993: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2994: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd2995: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2996: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd2997: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd2998: out = 32'b11010010100000000000000010000001; // MOVZ X1, 4
         16'd2999: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3000: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd3001: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3002: out = 32'b11110010100000101000101100000001; // MOVK X1, 5208
         16'd3003: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3004: out = 32'b11110010100010110000101100000001; // MOVK X1, 22616
         16'd3005: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3006: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3007: out = 32'b11010010100010110000000010000001; // MOVZ X1, 22532
         16'd3008: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3009: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3010: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3011: out = 32'b11110010100000000000100000000001; // MOVK X1, 64
         16'd3012: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3013: out = 32'b11110010100100101000100000000001; // MOVK X1, 37952
         16'd3014: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3015: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3016: out = 32'b11010010100010000000100000000001; // MOVZ X1, 16448
         16'd3017: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3018: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd3019: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3020: out = 32'b11110010100010100001001010000001; // MOVK X1, 20628
         16'd3021: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3022: out = 32'b11110010100100100001001000000001; // MOVK X1, 37008
         16'd3023: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3024: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3025: out = 32'b11010010100100100001001010000001; // MOVZ X1, 37012
         16'd3026: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3027: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd3028: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3029: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd3030: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3031: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd3032: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3033: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3034: out = 32'b11010010100111010001110100000001; // MOVZ X1, 59624
         16'd3035: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3036: out = 32'b11110010100111001001110010000001; // MOVK X1, 58596
         16'd3037: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3038: out = 32'b11110010100100101000101000000001; // MOVK X1, 37968
         16'd3039: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3040: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3041: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3042: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3043: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd3044: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3045: out = 32'b11110010100010100000100000000001; // MOVK X1, 20544
         16'd3046: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3047: out = 32'b11110010100000000000001000000001; // MOVK X1, 16
         16'd3048: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3049: out = 32'b11110010100000100000001000000001; // MOVK X1, 4112
         16'd3050: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3051: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3052: out = 32'b11010010100000100000101000000001; // MOVZ X1, 4176
         16'd3053: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3054: out = 32'b11110010100010100000101000000001; // MOVK X1, 20560
         16'd3055: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3056: out = 32'b11110010100010100000101010000001; // MOVK X1, 20564
         16'd3057: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3058: out = 32'b11110010100011001001010010000001; // MOVK X1, 25764
         16'd3059: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3060: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3061: out = 32'b11010010100101001001010100000001; // MOVZ X1, 42152
         16'd3062: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3063: out = 32'b11110010100101010000101010000001; // MOVK X1, 43092
         16'd3064: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3065: out = 32'b11110010100010100001011100000001; // MOVK X1, 20664
         16'd3066: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3067: out = 32'b11110010100101010000101000000001; // MOVK X1, 43088
         16'd3068: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3069: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3070: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3071: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3072: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3073: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3074: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd3075: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3076: out = 32'b11110010100010101000101100000001; // MOVK X1, 21592
         16'd3077: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3078: out = 32'b11110010100010110000101100000001; // MOVK X1, 22616
         16'd3079: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3080: out = 32'b11110010100010110000101100000001; // MOVK X1, 22616
         16'd3081: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3082: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3083: out = 32'b11010010100000001000000000000001; // MOVZ X1, 1024
         16'd3084: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3085: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3086: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3087: out = 32'b11110010100000000000100000000001; // MOVK X1, 64
         16'd3088: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3089: out = 32'b11110010100100100000100000000001; // MOVK X1, 36928
         16'd3090: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3091: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3092: out = 32'b11010010100010000000100000000001; // MOVZ X1, 16448
         16'd3093: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3094: out = 32'b11110010100000000000100000000001; // MOVK X1, 64
         16'd3095: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3096: out = 32'b11110010100010000001001010000001; // MOVK X1, 16532
         16'd3097: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3098: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd3099: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3100: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3101: out = 32'b11010010100100101001001010000001; // MOVZ X1, 38036
         16'd3102: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3103: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd3104: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3105: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd3106: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3107: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd3108: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3109: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3110: out = 32'b11010010100111010001110100000001; // MOVZ X1, 59624
         16'd3111: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3112: out = 32'b11110010100101001001001010000001; // MOVK X1, 42132
         16'd3113: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3114: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd3115: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3116: out = 32'b11110010100010100000101000000001; // MOVK X1, 20560
         16'd3117: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3118: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3119: out = 32'b11010010100010100000101010000001; // MOVZ X1, 20564
         16'd3120: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3121: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd3122: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3123: out = 32'b11110010100010100000000000000001; // MOVK X1, 20480
         16'd3124: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3125: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3126: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3127: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3128: out = 32'b11010010100010000000101000000001; // MOVZ X1, 16464
         16'd3129: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3130: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd3131: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3132: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3133: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3134: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3135: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3136: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3137: out = 32'b11010010100010100000100000000001; // MOVZ X1, 20544
         16'd3138: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3139: out = 32'b11110010100000000000101010000001; // MOVK X1, 84
         16'd3140: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3141: out = 32'b11110010100011001001011100000001; // MOVK X1, 25784
         16'd3142: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3143: out = 32'b11110010100111110001010010000001; // MOVK X1, 63652
         16'd3144: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3145: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3146: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3147: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3148: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3149: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3150: out = 32'b11010010100010101000000010000001; // MOVZ X1, 21508
         16'd3151: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3152: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd3153: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3154: out = 32'b11110010100010101000101100000001; // MOVK X1, 21592
         16'd3155: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3156: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd3157: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3158: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3159: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd3160: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3161: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3162: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3163: out = 32'b11110010100000000000100000000001; // MOVK X1, 64
         16'd3164: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3165: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd3166: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3167: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3168: out = 32'b11010010100010000000000000000001; // MOVZ X1, 16384
         16'd3169: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3170: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3171: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3172: out = 32'b11110010100010000001001010000001; // MOVK X1, 16532
         16'd3173: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3174: out = 32'b11110010100101001001110010000001; // MOVK X1, 42212
         16'd3175: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3176: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3177: out = 32'b11010010100111001001001010000001; // MOVZ X1, 58516
         16'd3178: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3179: out = 32'b11110010100100101001110010000001; // MOVK X1, 38116
         16'd3180: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3181: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd3182: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3183: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd3184: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3185: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3186: out = 32'b11010010100111010001010010000001; // MOVZ X1, 59556
         16'd3187: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3188: out = 32'b11110010100100101001010100000001; // MOVK X1, 38056
         16'd3189: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3190: out = 32'b11110010100111111001111110000001; // MOVK X1, 64764
         16'd3191: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3192: out = 32'b11110010100111111001111110000001; // MOVK X1, 64764
         16'd3193: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3194: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3195: out = 32'b11010010100111111001111110000001; // MOVZ X1, 64764
         16'd3196: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3197: out = 32'b11110010100111111001111110000001; // MOVK X1, 64764
         16'd3198: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3199: out = 32'b11110010100111111001111100000001; // MOVK X1, 64760
         16'd3200: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3201: out = 32'b11110010100101110001010100000001; // MOVK X1, 47272
         16'd3202: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3203: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3204: out = 32'b11010010100111010001110100000001; // MOVZ X1, 59624
         16'd3205: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3206: out = 32'b11110010100111010001010100000001; // MOVK X1, 59560
         16'd3207: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3208: out = 32'b11110010100101010000110010000001; // MOVK X1, 43108
         16'd3209: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3210: out = 32'b11110010100010101001010010000001; // MOVK X1, 21668
         16'd3211: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3212: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3213: out = 32'b11010010100111001001001010000001; // MOVZ X1, 58516
         16'd3214: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3215: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd3216: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3217: out = 32'b11110010100101001001010010000001; // MOVK X1, 42148
         16'd3218: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3219: out = 32'b11110010100101001001110100000001; // MOVK X1, 42216
         16'd3220: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3221: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3222: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3223: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3224: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3225: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3226: out = 32'b11010010100000001000000000000001; // MOVZ X1, 1024
         16'd3227: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3228: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3229: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3230: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3231: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3232: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3233: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3234: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3235: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd3236: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3237: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3238: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3239: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3240: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3241: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd3242: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3243: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3244: out = 32'b11010010100010000000100000000001; // MOVZ X1, 16448
         16'd3245: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3246: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3247: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3248: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd3249: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3250: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd3251: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3252: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3253: out = 32'b11010010100111001001110100000001; // MOVZ X1, 58600
         16'd3254: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3255: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd3256: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3257: out = 32'b11110010100111010001111100000001; // MOVK X1, 59640
         16'd3258: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3259: out = 32'b11110010100111110001110100000001; // MOVK X1, 63720
         16'd3260: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3261: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3262: out = 32'b11010010100100101001001010000001; // MOVZ X1, 38036
         16'd3263: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3264: out = 32'b11110010100100101001111110000001; // MOVK X1, 38140
         16'd3265: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3266: out = 32'b11110010100111111001111110000001; // MOVK X1, 64764
         16'd3267: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3268: out = 32'b11110010100111111001111110000001; // MOVK X1, 64764
         16'd3269: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3270: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3271: out = 32'b11111000000000000000000001001110; // STUR X14, [X2, 0]
         16'd3272: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3273: out = 32'b11111000000000000000000001001110; // STUR X14, [X2, 0]
         16'd3274: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3275: out = 32'b11111000000000000000000001001110; // STUR X14, [X2, 0]
         16'd3276: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3277: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3278: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3279: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3280: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3281: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3282: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3283: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd3284: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3285: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3286: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3287: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3288: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3289: out = 32'b11110010100000000000100000000001; // MOVK X1, 64
         16'd3290: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3291: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3292: out = 32'b11010010100010000000100000000001; // MOVZ X1, 16448
         16'd3293: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3294: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3295: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3296: out = 32'b11110010100000000000100000000001; // MOVK X1, 64
         16'd3297: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3298: out = 32'b11110010100010000001001010000001; // MOVK X1, 16532
         16'd3299: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3300: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3301: out = 32'b11010010100100101001110010000001; // MOVZ X1, 38116
         16'd3302: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3303: out = 32'b11110010100111001001110100000001; // MOVK X1, 58600
         16'd3304: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3305: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd3306: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3307: out = 32'b11110010100111010001010010000001; // MOVK X1, 59556
         16'd3308: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3309: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3310: out = 32'b11010010100100101000101010000001; // MOVZ X1, 37972
         16'd3311: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3312: out = 32'b11110010100010101000110100000001; // MOVK X1, 21608
         16'd3313: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3314: out = 32'b11110010100011010001010110000001; // MOVK X1, 26796
         16'd3315: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3316: out = 32'b11110010100101011001010110000001; // MOVK X1, 44204
         16'd3317: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3318: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3319: out = 32'b11010010100101111001011110000001; // MOVZ X1, 48316
         16'd3320: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3321: out = 32'b11110010100101111001011110000001; // MOVK X1, 48316
         16'd3322: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3323: out = 32'b11110010100101111001011110000001; // MOVK X1, 48316
         16'd3324: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3325: out = 32'b11110010100111111001111110000001; // MOVK X1, 64764
         16'd3326: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3327: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3328: out = 32'b11111000000000000000000001001110; // STUR X14, [X2, 0]
         16'd3329: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3330: out = 32'b11111000000000000000000001001110; // STUR X14, [X2, 0]
         16'd3331: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3332: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3333: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3334: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3335: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3336: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3337: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3338: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3339: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3340: out = 32'b11010010100000000000100000000001; // MOVZ X1, 64
         16'd3341: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3342: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3343: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3344: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3345: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3346: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd3347: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3348: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3349: out = 32'b11010010100100101001001010000001; // MOVZ X1, 38036
         16'd3350: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3351: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd3352: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3353: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd3354: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3355: out = 32'b11110010100101001001001010000001; // MOVK X1, 42132
         16'd3356: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3357: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3358: out = 32'b11010010100010100000101000000001; // MOVZ X1, 20560
         16'd3359: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3360: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3361: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3362: out = 32'b11110010100000000000000010000001; // MOVK X1, 4
         16'd3363: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3364: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd3365: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3366: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3367: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd3368: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3369: out = 32'b11110010100000101000001010000001; // MOVK X1, 5140
         16'd3370: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3371: out = 32'b11110010100000101000101010000001; // MOVK X1, 5204
         16'd3372: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3373: out = 32'b11110010100010101000101010000001; // MOVK X1, 21588
         16'd3374: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3375: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3376: out = 32'b11010010100010110000101100000001; // MOVZ X1, 22616
         16'd3377: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3378: out = 32'b11110010100010110000110100000001; // MOVK X1, 22632
         16'd3379: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3380: out = 32'b11110010100011010001010100000001; // MOVK X1, 26792
         16'd3381: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3382: out = 32'b11110010100101010001010100000001; // MOVK X1, 43176
         16'd3383: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3384: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3385: out = 32'b11010010100101011001010110000001; // MOVZ X1, 44204
         16'd3386: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3387: out = 32'b11110010100101011001011110000001; // MOVK X1, 44220
         16'd3388: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3389: out = 32'b11110010100101111001011110000001; // MOVK X1, 48316
         16'd3390: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3391: out = 32'b11110010100101111001011110000001; // MOVK X1, 48316
         16'd3392: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3393: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3394: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3395: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3396: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3397: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3398: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3399: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3400: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3401: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3402: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3403: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3404: out = 32'b11010010100010000000100000000001; // MOVZ X1, 16448
         16'd3405: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3406: out = 32'b11110010100010000000101010000001; // MOVK X1, 16468
         16'd3407: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3408: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd3409: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3410: out = 32'b11110010100010100000101000000001; // MOVK X1, 20560
         16'd3411: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3412: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3413: out = 32'b11010010100100101000100000000001; // MOVZ X1, 37952
         16'd3414: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3415: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3416: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3417: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3418: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3419: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3420: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3421: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3422: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3423: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3424: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd3425: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3426: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd3427: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3428: out = 32'b11110010100000000000000010000001; // MOVK X1, 4
         16'd3429: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3430: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd3431: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3432: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3433: out = 32'b11010010100000001000000000000001; // MOVZ X1, 1024
         16'd3434: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3435: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3436: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3437: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd3438: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3439: out = 32'b11110010100000001000001010000001; // MOVK X1, 1044
         16'd3440: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3441: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3442: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3443: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3444: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3445: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3446: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3447: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3448: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3449: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3450: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3451: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3452: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd3453: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3454: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3455: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3456: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd3457: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3458: out = 32'b11110010100010100001001010000001; // MOVK X1, 20628
         16'd3459: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3460: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3461: out = 32'b11010010100100101000000000000001; // MOVZ X1, 37888
         16'd3462: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3463: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3464: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3465: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3466: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3467: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3468: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3469: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3470: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3471: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3472: out = 32'b11010010100000001000000010000001; // MOVZ X1, 1028
         16'd3473: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3474: out = 32'b11110010100000001000000000000001; // MOVK X1, 1024
         16'd3475: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3476: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3477: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3478: out = 32'b11110010100000001000000010000001; // MOVK X1, 1028
         16'd3479: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3480: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3481: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3482: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3483: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3484: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3485: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3486: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3487: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3488: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3489: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3490: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3491: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3492: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3493: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd3494: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3495: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3496: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3497: out = 32'b11110010100000000000101000000001; // MOVK X1, 80
         16'd3498: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3499: out = 32'b11110010100100101001110100000001; // MOVK X1, 38120
         16'd3500: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3501: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3502: out = 32'b11010010100010101000000000000001; // MOVZ X1, 21504
         16'd3503: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3504: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3505: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3506: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3507: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3508: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3509: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3510: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3511: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3512: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3513: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3514: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3515: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3516: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3517: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3518: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3519: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3520: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3521: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3522: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3523: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3524: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3525: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3526: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3527: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd3528: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3529: out = 32'b11110010100000000000100000000001; // MOVK X1, 64
         16'd3530: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3531: out = 32'b11110010100010100001001010000001; // MOVK X1, 20628
         16'd3532: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3533: out = 32'b11110010100111001001010100000001; // MOVK X1, 58536
         16'd3534: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3535: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3536: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3537: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3538: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3539: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3540: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3541: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3542: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3543: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3544: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3545: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3546: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3547: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3548: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3549: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3550: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3551: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3552: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3553: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3554: out = 32'b11010010100000000000100000000001; // MOVZ X1, 64
         16'd3555: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3556: out = 32'b11110010100010101001001010000001; // MOVK X1, 21652
         16'd3557: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3558: out = 32'b11110010100101001001110010000001; // MOVK X1, 42212
         16'd3559: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3560: out = 32'b11110010100111010001010010000001; // MOVK X1, 59556
         16'd3561: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3562: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3563: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd3564: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3565: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3566: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3567: out = 32'b11110010100010000000000000000001; // MOVK X1, 16384
         16'd3568: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3569: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3570: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3571: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3572: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3573: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3574: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3575: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3576: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3577: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3578: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3579: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3580: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3581: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3582: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3583: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3584: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3585: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3586: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd3587: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3588: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3589: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3590: out = 32'b11110010100000000000100000000001; // MOVK X1, 64
         16'd3591: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3592: out = 32'b11110010100010000000100000000001; // MOVK X1, 16448
         16'd3593: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3594: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3595: out = 32'b11010010100010101001001010000001; // MOVZ X1, 21652
         16'd3596: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3597: out = 32'b11110010100101001001010010000001; // MOVK X1, 42148
         16'd3598: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3599: out = 32'b11110010100101001001110010000001; // MOVK X1, 42212
         16'd3600: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3601: out = 32'b11110010100111010000101010000001; // MOVK X1, 59476
         16'd3602: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3603: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3604: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd3605: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3606: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3607: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3608: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3609: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3610: out = 32'b11110010100010000000000000000001; // MOVK X1, 16384
         16'd3611: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3612: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3613: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3614: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3615: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3616: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3617: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3618: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3619: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3620: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3621: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3622: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3623: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3624: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3625: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3626: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3627: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd3628: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3629: out = 32'b11110010100000000000100000000001; // MOVK X1, 64
         16'd3630: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3631: out = 32'b11110010100010101001001010000001; // MOVK X1, 21652
         16'd3632: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3633: out = 32'b11110010100100101001001010000001; // MOVK X1, 38036
         16'd3634: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3635: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3636: out = 32'b11010010100010100001001010000001; // MOVZ X1, 20628
         16'd3637: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3638: out = 32'b11110010100101001001010010000001; // MOVK X1, 42148
         16'd3639: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3640: out = 32'b11110010100111001001110100000001; // MOVK X1, 58600
         16'd3641: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3642: out = 32'b11110010100111010000101000000001; // MOVK X1, 59472
         16'd3643: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3644: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3645: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3646: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3647: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3648: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3649: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3650: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3651: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3652: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3653: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3654: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3655: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3656: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3657: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3658: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3659: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3660: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3661: out = 32'b11010010100000000000100000000001; // MOVZ X1, 64
         16'd3662: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3663: out = 32'b11110010100100101001010010000001; // MOVK X1, 38052
         16'd3664: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3665: out = 32'b11110010100101010001010010000001; // MOVK X1, 43172
         16'd3666: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3667: out = 32'b11110010100101001001001010000001; // MOVK X1, 42132
         16'd3668: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3669: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3670: out = 32'b11010010100010100001001010000001; // MOVZ X1, 20628
         16'd3671: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3672: out = 32'b11110010100100101001010010000001; // MOVK X1, 38052
         16'd3673: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3674: out = 32'b11110010100111001001110100000001; // MOVK X1, 58600
         16'd3675: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3676: out = 32'b11110010100101010000100000000001; // MOVK X1, 43072
         16'd3677: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3678: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3679: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3680: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3681: out = 32'b11010010100010000000000000000001; // MOVZ X1, 16384
         16'd3682: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3683: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3684: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3685: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3686: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3687: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3688: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3689: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3690: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3691: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3692: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3693: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3694: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3695: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3696: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3697: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3698: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3699: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3700: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3701: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3702: out = 32'b11010010100100101001010010000001; // MOVZ X1, 38052
         16'd3703: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3704: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd3705: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3706: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd3707: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3708: out = 32'b11110010100101001001001010000001; // MOVK X1, 42132
         16'd3709: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3710: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3711: out = 32'b11010010100100101001001010000001; // MOVZ X1, 38036
         16'd3712: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3713: out = 32'b11110010100100101001010010000001; // MOVK X1, 38052
         16'd3714: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3715: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd3716: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3717: out = 32'b11110010100100101000000000000001; // MOVK X1, 37888
         16'd3718: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3719: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3720: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3721: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3722: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3723: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3724: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3725: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3726: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3727: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3728: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3729: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3730: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3731: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3732: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3733: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3734: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3735: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3736: out = 32'b11010010100100101001110100000001; // MOVZ X1, 38120
         16'd3737: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3738: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd3739: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3740: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd3741: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3742: out = 32'b11110010100111010001010010000001; // MOVK X1, 59556
         16'd3743: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3744: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3745: out = 32'b11010010100100101001001010000001; // MOVZ X1, 38036
         16'd3746: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3747: out = 32'b11110010100101001001110100000001; // MOVK X1, 42216
         16'd3748: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3749: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd3750: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3751: out = 32'b11110010100010101000000000000001; // MOVK X1, 21504
         16'd3752: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3753: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3754: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3755: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3756: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3757: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3758: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3759: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3760: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3761: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3762: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3763: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3764: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3765: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3766: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3767: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3768: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3769: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3770: out = 32'b11010010100000000001001010000001; // MOVZ X1, 148
         16'd3771: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3772: out = 32'b11110010100111110001110100000001; // MOVK X1, 63720
         16'd3773: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3774: out = 32'b11110010100111010001110100000001; // MOVK X1, 59624
         16'd3775: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3776: out = 32'b11110010100111010001010010000001; // MOVK X1, 59556
         16'd3777: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3778: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3779: out = 32'b11010010100101001001010010000001; // MOVZ X1, 42148
         16'd3780: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3781: out = 32'b11110010100111001001110100000001; // MOVK X1, 58600
         16'd3782: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3783: out = 32'b11110010100111010001010100000001; // MOVK X1, 59560
         16'd3784: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3785: out = 32'b11110010100010000000000000000001; // MOVK X1, 16384
         16'd3786: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3787: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3788: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3789: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3790: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3791: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3792: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3793: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3794: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd3795: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3796: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3797: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3798: out = 32'b11110010100000000000100000000001; // MOVK X1, 64
         16'd3799: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3800: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3801: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3802: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3803: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3804: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3805: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3806: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3807: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3808: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3809: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3810: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3811: out = 32'b11010010100000000000000000000001; // MOVZ X1, 0
         16'd3812: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3813: out = 32'b11110010100100101001111100000001; // MOVK X1, 38136
         16'd3814: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3815: out = 32'b11110010100111110001111100000001; // MOVK X1, 63736
         16'd3816: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3817: out = 32'b11110010100111010001010010000001; // MOVK X1, 59556
         16'd3818: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3819: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3820: out = 32'b11010010100101001001010010000001; // MOVZ X1, 42148
         16'd3821: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3822: out = 32'b11110010100111001001110100000001; // MOVK X1, 58600
         16'd3823: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3824: out = 32'b11110010100111010001001010000001; // MOVK X1, 59540
         16'd3825: out = 32'b11010011011000000100000000100001; // LSL X1, X1, 16
         16'd3826: out = 32'b11110010100000000000000000000001; // MOVK X1, 0
         16'd3827: out = 32'b11111000000000000000000001000001; // STUR X1, [X2, 0]
         16'd3828: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3829: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3830: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3831: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3832: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3833: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3834: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3835: out = 32'b11111000000000000000000001010010; // STUR X18, [X2, 0]
         16'd3836: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
         16'd3837: out = 32'b11010010100000000000000010100101; // MOVZ X5, 5
         16'd3838: out = 32'b11111000000000000000001010000101; // STUR X5, [X20, 0]
         16'd3839: out = 32'b00010111111111111111111111111111; // B -1
         default: out = 32'b11010110000000000000001111100000; // BR XZR
      endcase
   end
endmodule
