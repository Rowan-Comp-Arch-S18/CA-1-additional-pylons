module KeyboardV3(CLOCK_50, PS2_KBCLK, PS2_KBDAT, REG0, REG1);
	input CLOCK_50;														// Board clock
   input PS2_KBCLK;														// Keyboard clock
   input PS2_KBDAT;														// Keyboard data
	
   output reg [63:0] REG0;
	output reg [63:0] REG1;
	
	reg CLOCK_DOWN250;													// CLOCK_50/250
	reg [6:0] CLOCK_COUNTER; 											// Counter for dividing CLOCK_50
	reg LAST_KBCLK;														// Stores last state of PS2_KBCLK
	reg [10:0] SCANNED_PACKET;											// Stores incoming packet
	reg [3:0] PACKET_COUNTER;											// Counts number of bits in the incoming packet
	reg [63:0] TIMEOUT_COUNTER;										// Counter for timeout
	reg TIMEOUT;															// True after 1/10 sec of no input
	
	parameter KB_ESC = 8'h76, KB_F1 = 8'h05, KB_F2 = 8'h06, 
	KB_F3 = 8'h04, KB_F4 = 8'h0C, KB_F5 = 8'h03, 
	KB_F6 = 8'h0B, KB_F7 = 8'h83, KB_F8 = 8'h0A, 
	KB_F9 = 8'h01, KB_F10 = 8'h09, KB_F11 = 8'h78, 
	KB_F12 = 8'h07, KB_GRAVE = 8'h0E, KB_1 = 8'h16, 
	KB_2 = 8'h1E, KB_3 = 8'h26, KB_4 = 8'h25, KB_5 = 8'h2E, 
	KB_6 = 8'h36, KB_7 = 8'h3D, KB_8 = 8'h3E, KB_9 = 8'h46, 
	KB_0 = 8'h45, KB_MINUS = 8'h4E, KB_EQUALS = 8'h55, 
	KB_BACKSPACE = 8'h66, KB_TAB = 8'h0D, KB_Q = 8'h15, 
	KB_W = 8'h1D, KB_E = 8'h24, KB_R = 8'h2D, KB_T = 8'h2C, 
	KB_Y = 8'h35, KB_U = 8'h3C, KB_I = 8'h43, KB_O = 9'h44, 
	KB_P = 8'h4D, KB_LEFTBRACKET = 8'h54, 
	KB_RIGHTBRACKET = 8'h5B, KB_BLACKSLASH = 8'h5D, 
	KB_CAPS = 8'h58, KB_A = 8'h1C, KB_S = 8'h1B, 
	KB_D = 8'h23, KB_F = 8'h2B, KB_G = 8'h34, KB_H = 8'h33, 
	KB_J = 8'h3B, KB_K = 8'h42, KB_L = 8'h4B, 
	KB_SEMICOLON = 8'h4C, KB_APOSTROPHE = 8'h52, 
	KB_ENTER = 8'h5A, KB_LEFTSHIFT = 8'h12, KB_Z = 8'h1A, 
	KB_X = 8'h22, KB_C = 8'h21, KB_V = 8'h2A, KB_B = 8'h32, 
	KB_N = 8'h31, KB_M = 8'h3A, KB_COMMA = 8'h41, 
	KB_PERIOD = 8'h49, KB_SLASH = 8'h4A, 
	KB_RIGHTSHIFT = 8'h59, KB_CTRL = 8'h14, KB_ALT = 8'h11, 
	KB_SPACE = 8'h29, KB_UP = 8'h75, KB_LEFT = 8'h6B, 
	KB_DOWN = 8'h72, KB_RIGHT = 8'h74;
	
	initial begin
		CLOCK_DOWN250 <= 1'd0;
		CLOCK_COUNTER <= 7'd0;
		LAST_KBCLK <= 1'd0;
		SCANNED_PACKET <= 11'd0;
		PACKET_COUNTER <= 4'd0;
		TIMEOUT_COUNTER <= 64'd0;
		TIMEOUT <= 1'd0;
		REG0 <= 64'd0;
		REG1 <= 64'd0;
	end
	
	always @(posedge CLOCK_50) begin
		if (CLOCK_COUNTER > 124) begin
			CLOCK_DOWN250 <= ~CLOCK_DOWN250;
			CLOCK_COUNTER <= 7'd0;
		end
		else begin
			CLOCK_COUNTER <= CLOCK_COUNTER + 1'd1;
		end
	end
	
	always @(posedge CLOCK_DOWN250) begin
		if (TIMEOUT_COUNTER > 20000)
			TIMEOUT <= 1'd1;
		else
			TIMEOUT <= 1'd0;
	end
	
	always @(posedge CLOCK_DOWN250) begin
		if (PS2_KBCLK != LAST_KBCLK) begin
			TIMEOUT_COUNTER <= 64'd0;
			if (PS2_KBCLK == 0) begin
				PACKET_COUNTER <= PACKET_COUNTER + 1'd1;
				SCANNED_PACKET <= {PS2_KBDAT, SCANNED_PACKET[10:1]};
			end
			else begin
				if (PACKET_COUNTER == 11) begin
					
					if (SCANNED_PACKET[8:1] == KB_ESC) begin
						REG0 <= 64'b0000000000000000000000000000000000000000000000000000000000000001;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_F1) begin
						REG0 <= 64'b0000000000000000000000000000000000000000000000000000000000000010;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_F2) begin
						REG0 <= 64'b0000000000000000000000000000000000000000000000000000000000000100;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_F3) begin
						REG0 <= 64'b0000000000000000000000000000000000000000000000000000000000001000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_F4) begin
						REG0 <= 64'b0000000000000000000000000000000000000000000000000000000000010000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_F5) begin
						REG0 <= 64'b0000000000000000000000000000000000000000000000000000000000100000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_F6) begin
						REG0 <= 64'b0000000000000000000000000000000000000000000000000000000001000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_F7) begin
						REG0 <= 64'b0000000000000000000000000000000000000000000000000000000010000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_F8) begin
						REG0 <= 64'b0000000000000000000000000000000000000000000000000000000100000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_F9) begin
						REG0 <= 64'b0000000000000000000000000000000000000000000000000000001000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_F10) begin
						REG0 <= 64'b0000000000000000000000000000000000000000000000000000010000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_F11) begin
						REG0 <= 64'b0000000000000000000000000000000000000000000000000000100000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_F12) begin
						REG0 <= 64'b0000000000000000000000000000000000000000000000000001000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_GRAVE) begin
						REG0 <= 64'b0000000000000000000000000000000000000000000000000010000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_1) begin
						REG0 <= 64'b0000000000000000000000000000000000000000000000000100000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_2) begin
						REG0 <= 64'b0000000000000000000000000000000000000000000000001000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_3) begin
						REG0 <= 64'b0000000000000000000000000000000000000000000000010000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_4) begin
						REG0 <= 64'b0000000000000000000000000000000000000000000000100000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_5) begin
						REG0 <= 64'b0000000000000000000000000000000000000000000001000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_6) begin
						REG0 <= 64'b0000000000000000000000000000000000000000000010000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_7) begin
						REG0 <= 64'b0000000000000000000000000000000000000000000100000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_8) begin
						REG0 <= 64'b0000000000000000000000000000000000000000001000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_9) begin
						REG0 <= 64'b0000000000000000000000000000000000000000010000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_0) begin
						REG0 <= 64'b0000000000000000000000000000000000000000100000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_MINUS) begin
						REG0 <= 64'b0000000000000000000000000000000000000001000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_EQUALS) begin
						REG0 <= 64'b0000000000000000000000000000000000000010000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_BACKSPACE) begin
						REG0 <= 64'b0000000000000000000000000000000000000100000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_TAB) begin
						REG0 <= 64'b0000000000000000000000000000000000001000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_Q) begin
						REG0 <= 64'b0000000000000000000000000000000000010000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_W) begin
						REG0 <= 64'b0000000000000000000000000000000000100000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_E) begin
						REG0 <= 64'b0000000000000000000000000000000001000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_R) begin
						REG0 <= 64'b0000000000000000000000000000000010000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_T) begin
						REG0 <= 64'b0000000000000000000000000000000100000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_Y) begin
						REG0 <= 64'b0000000000000000000000000000001000000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_U) begin
						REG0 <= 64'b0000000000000000000000000000010000000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_I) begin
						REG0 <= 64'b0000000000000000000000000000100000000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_O) begin
						REG0 <= 64'b0000000000000000000000000001000000000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_P) begin
						REG0 <= 64'b0000000000000000000000000010000000000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_LEFTBRACKET) begin
						REG0 <= 64'b0000000000000000000000000100000000000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_RIGHTBRACKET) begin
						REG0 <= 64'b0000000000000000000000001000000000000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_BLACKSLASH) begin
						REG0 <= 64'b0000000000000000000000010000000000000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_CAPS) begin
						REG0 <= 64'b0000000000000000000000100000000000000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_A) begin
						REG0 <= 64'b0000000000000000000001000000000000000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_S) begin
						REG0 <= 64'b0000000000000000000010000000000000000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_D) begin
						REG0 <= 64'b0000000000000000000100000000000000000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_F) begin
						REG0 <= 64'b0000000000000000001000000000000000000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_G) begin
						REG0 <= 64'b0000000000000000010000000000000000000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_H) begin
						REG0 <= 64'b0000000000000000100000000000000000000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_J) begin
						REG0 <= 64'b0000000000000001000000000000000000000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_K) begin
						REG0 <= 64'b0000000000000010000000000000000000000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_L) begin
						REG0 <= 64'b0000000000000100000000000000000000000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_SEMICOLON) begin
						REG0 <= 64'b0000000000001000000000000000000000000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_APOSTROPHE) begin
						REG0 <= 64'b0000000000010000000000000000000000000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_ENTER) begin
						REG0 <= 64'b0000000000100000000000000000000000000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_LEFTSHIFT) begin
						REG0 <= 64'b0000000001000000000000000000000000000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_Z) begin
						REG0 <= 64'b0000000010000000000000000000000000000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_X) begin
						REG0 <= 64'b0000000100000000000000000000000000000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_C) begin
						REG0 <= 64'b0000001000000000000000000000000000000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_V) begin
						REG0 <= 64'b0000010000000000000000000000000000000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_B) begin
						REG0 <= 64'b0000100000000000000000000000000000000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_N) begin
						REG0 <= 64'b0001000000000000000000000000000000000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_M) begin
						REG0 <= 64'b0010000000000000000000000000000000000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_COMMA) begin
						REG0 <= 64'b0100000000000000000000000000000000000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_PERIOD) begin
						REG0 <= 64'b1000000000000000000000000000000000000000000000000000000000000000;
						REG1 <= 64'd0;
					end
					else if (SCANNED_PACKET[8:1] == KB_SLASH) begin
						REG0 <= 64'd0;
						REG1 <= 64'b0000000000000000000000000000000000000000000000000000000000000001;
					end
					else if (SCANNED_PACKET[8:1] == KB_RIGHTSHIFT) begin
						REG0 <= 64'd0;
						REG1 <= 64'b0000000000000000000000000000000000000000000000000000000000000010;
					end
					else if (SCANNED_PACKET[8:1] == KB_CTRL) begin
						REG0 <= 64'd0;
						REG1 <= 64'b0000000000000000000000000000000000000000000000000000000000000100;
					end
					else if (SCANNED_PACKET[8:1] == KB_ALT) begin
						REG0 <= 64'd0;
						REG1 <= 64'b0000000000000000000000000000000000000000000000000000000000001000;
					end
					else if (SCANNED_PACKET[8:1] == KB_SPACE) begin
						REG0 <= 64'd0;
						REG1 <= 64'b0000000000000000000000000000000000000000000000000000000000010000;
					end
					else if (SCANNED_PACKET[8:1] == KB_UP) begin
						REG0 <= 64'd0;
						REG1 <= 64'b0000000000000000000000000000000000000000000000000000000000100000;
					end
					else if (SCANNED_PACKET[8:1] == KB_LEFT) begin
						REG0 <= 64'd0;
						REG1 <= 64'b0000000000000000000000000000000000000000000000000000000001000000;
					end
					else if (SCANNED_PACKET[8:1] == KB_DOWN) begin
						REG0 <= 64'd0;
						REG1 <= 64'b0000000000000000000000000000000000000000000000000000000010000000;
					end
					else if (SCANNED_PACKET[8:1] == KB_RIGHT) begin
						REG0 <= 64'd0;
						REG1 <= 64'b0000000000000000000000000000000000000000000000000000000100000000;
					end
					
					PACKET_COUNTER <= 0;
				end
			end
		end
		if (PS2_KBCLK == LAST_KBCLK) begin
			TIMEOUT_COUNTER <= TIMEOUT_COUNTER + 1'd1;
			if (TIMEOUT) begin
				REG0 <= 64'd0;
				REG1 <= 64'd0;
				PACKET_COUNTER <= 0;
				TIMEOUT_COUNTER <= 64'd0;
			end
		end
		LAST_KBCLK <= PS2_KBCLK;
	end
endmodule
