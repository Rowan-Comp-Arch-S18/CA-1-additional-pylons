module GPUCharDecoder(row, col, char, charPixelOn);
	input [3:0] row;
	input [2:0] col;
	input [7:0] char;
	output charPixelOn;
	
	// TODO
	assign charPixelOn = 1'b1;
endmodule
