module InstructionReg();